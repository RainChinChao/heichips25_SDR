module heichips25_template (clk,
    ena,
    rst_n,
    VPWR,
    VGND,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 inout VPWR;
 inout VGND;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire \Demo1.epsk_de1.bit_out[0] ;
 wire \Demo1.epsk_de1.bit_out[1] ;
 wire \Demo1.epsk_de1.bit_out[2] ;
 wire \Demo1.qam16_bits[0] ;
 wire \Demo1.qam16_bits[1] ;
 wire \Demo1.qam16_bits[2] ;
 wire \Demo1.qam16_bits[3] ;
 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire net38;
 wire \mod1.bpsk_mod.i_out[2] ;
 wire \mod1.i_out_8psk[0] ;
 wire \mod1.i_out_8psk[1] ;
 wire \mod1.i_out_8psk[2] ;
 wire \mod1.i_out_qam16[2] ;
 wire \mod1.i_out_qam16[3] ;
 wire \mod1.i_out_qpsk[1] ;
 wire \mod1.i_out_qpsk[2] ;
 wire \mod1.psk8_mod.q_out[1] ;
 wire \mod1.psk8_mod.q_out[2] ;
 wire \mod1.q_out_qam16[2] ;
 wire \mod1.q_out_qam16[3] ;
 wire \mod1.q_out_qpsk[2] ;
 wire \mod1.qam16_mod.i_level[2] ;
 wire \mod1.qam16_mod.i_level[3] ;
 wire \mod1.qam16_mod.q_level[2] ;
 wire \mod1.qam16_mod.q_level[3] ;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire clknet_0_clk;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net33;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire net46;
 wire net47;
 wire net48;

 sg13g2_inv_1 _055_ (.VDD(VPWR),
    .Y(\mod1.qam16_mod.q_level[3] ),
    .A(net3),
    .VSS(VGND));
 sg13g2_inv_1 _056_ (.VDD(VPWR),
    .Y(_032_),
    .A(net4),
    .VSS(VGND));
 sg13g2_inv_4 _057_ (.A(net5),
    .Y(\mod1.qam16_mod.i_level[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _058_ (.VDD(VPWR),
    .Y(_033_),
    .A(net7),
    .VSS(VGND));
 sg13g2_inv_1 _059_ (.VDD(VPWR),
    .Y(_034_),
    .A(net6),
    .VSS(VGND));
 sg13g2_inv_1 _060_ (.VDD(VPWR),
    .Y(_035_),
    .A(net47),
    .VSS(VGND));
 sg13g2_and2_1 _061_ (.A(net7),
    .B(net6),
    .X(_036_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _062_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_037_),
    .B(net10),
    .A(net16));
 sg13g2_and2_1 _063_ (.A(net9),
    .B(net8),
    .X(_038_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _064_ (.B1(net12),
    .VDD(VPWR),
    .Y(_011_),
    .VSS(VGND),
    .A1(_037_),
    .A2(_038_));
 sg13g2_nand2_2 _065_ (.Y(_039_),
    .A(_032_),
    .B(\mod1.qam16_mod.i_level[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _066_ (.A(net3),
    .B(net4),
    .Y(_040_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3b_1 _067_ (.B(\mod1.qam16_mod.i_level[3] ),
    .C(_040_),
    .Y(_000_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(net2));
 sg13g2_nor2b_2 _068_ (.A(net6),
    .B_N(net7),
    .Y(_041_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _069_ (.Y(_042_),
    .B1(_041_),
    .B2(\Demo1.epsk_de1.bit_out[0] ),
    .A2(net11),
    .A1(\Demo1.qam16_bits[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 _070_ (.A(_042_),
    .Y(net21),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _071_ (.Y(_043_),
    .B1(_041_),
    .B2(\Demo1.epsk_de1.bit_out[1] ),
    .A2(net11),
    .A1(\Demo1.qam16_bits[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 _072_ (.A(_043_),
    .Y(net22),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _073_ (.Y(_044_),
    .B1(_041_),
    .B2(\Demo1.epsk_de1.bit_out[2] ),
    .A2(net12),
    .A1(\Demo1.qam16_bits[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _074_ (.Y(net23),
    .A(_044_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _075_ (.A(\Demo1.qam16_bits[3] ),
    .B(net11),
    .X(net24),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _076_ (.B(net5),
    .A(net4),
    .X(\mod1.qam16_mod.i_level[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _077_ (.A(\mod1.i_out_8psk[0] ),
    .B(_041_),
    .X(net29),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _078_ (.A(net7),
    .B_N(net6),
    .Y(_045_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _079_ (.Y(_046_),
    .B1(_045_),
    .B2(\mod1.i_out_qpsk[1] ),
    .A2(net11),
    .A1(\Demo1.qam16_bits[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _080_ (.B1(_034_),
    .VDD(VPWR),
    .Y(_047_),
    .VSS(VGND),
    .A1(_033_),
    .A2(\mod1.i_out_8psk[1] ));
 sg13g2_nor3_1 _081_ (.A(net7),
    .B(net6),
    .C(\Demo1.qam16_bits[3] ),
    .Y(_048_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _082_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_048_),
    .Y(net26),
    .A2(_047_),
    .A1(_046_));
 sg13g2_nand2_1 _083_ (.Y(_049_),
    .A(\mod1.i_out_8psk[2] ),
    .B(_041_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _084_ (.Y(_050_),
    .A(\mod1.i_out_qpsk[2] ),
    .B(_045_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _085_ (.B(_034_),
    .C(\mod1.bpsk_mod.i_out[2] ),
    .A(_033_),
    .Y(_051_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _086_ (.Y(_052_),
    .A(\mod1.i_out_qam16[2] ),
    .B(net11),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _087_ (.B(_050_),
    .C(_051_),
    .A(_049_),
    .Y(net27),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_052_));
 sg13g2_nand2_1 _088_ (.Y(_053_),
    .A(\mod1.i_out_qam16[3] ),
    .B(net11),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _089_ (.B(_050_),
    .C(_051_),
    .A(_049_),
    .Y(net28),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_053_));
 sg13g2_nand2_1 _090_ (.Y(_015_),
    .A(\mod1.psk8_mod.q_out[1] ),
    .B(_041_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _091_ (.Y(net30),
    .A(_046_),
    .B(_015_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _092_ (.Y(_016_),
    .B1(_045_),
    .B2(\mod1.q_out_qpsk[2] ),
    .A2(_041_),
    .A1(\mod1.psk8_mod.q_out[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _093_ (.Y(_017_),
    .A(\mod1.q_out_qam16[2] ),
    .B(net11),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _094_ (.Y(net31),
    .A(_016_),
    .B(_017_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _095_ (.Y(_018_),
    .A(\mod1.q_out_qam16[3] ),
    .B(net11),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _096_ (.Y(net32),
    .A(_016_),
    .B(_018_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _097_ (.A(\mod1.qam16_mod.q_level[3] ),
    .B(net2),
    .Y(_019_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _098_ (.Y(_020_),
    .B(net3),
    .A_N(net2),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _099_ (.B(net2),
    .A(net3),
    .X(\mod1.qam16_mod.q_level[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _100_ (.Y(_021_),
    .A(net4),
    .B(\mod1.qam16_mod.q_level[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _101_ (.A(net5),
    .B(_021_),
    .Y(_006_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _102_ (.B(net4),
    .C(\mod1.qam16_mod.i_level[3] ),
    .A(net3),
    .Y(_022_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _103_ (.B1(_022_),
    .VDD(VPWR),
    .Y(_007_),
    .VSS(VGND),
    .A1(net2),
    .A2(_039_));
 sg13g2_o21ai_1 _104_ (.B1(_022_),
    .VDD(VPWR),
    .Y(_008_),
    .VSS(VGND),
    .A1(_039_),
    .A2(_020_));
 sg13g2_nor3_1 _105_ (.A(net5),
    .B(_040_),
    .C(_019_),
    .Y(_009_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _106_ (.A(_032_),
    .B(net5),
    .C(_019_),
    .Y(_010_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _107_ (.A(net20),
    .B(net12),
    .X(_023_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _108_ (.VDD(VPWR),
    .Y(_005_),
    .A(_023_),
    .VSS(VGND));
 sg13g2_or2_1 _109_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_024_),
    .B(net1),
    .A(net17));
 sg13g2_nand3_1 _110_ (.B(net18),
    .C(_024_),
    .A(net19),
    .Y(_025_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _111_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_026_),
    .B(net18),
    .A(net19));
 sg13g2_a21o_1 _112_ (.A2(net1),
    .A1(net17),
    .B1(_026_),
    .X(_027_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _113_ (.A(net20),
    .B_N(net12),
    .Y(_028_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _114_ (.Y(_004_),
    .B1(_027_),
    .B2(_028_),
    .A2(_025_),
    .A1(_023_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _115_ (.A(net19),
    .B(net18),
    .C(net17),
    .D(net1),
    .Y(_029_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _116_ (.A(_033_),
    .B(net6),
    .C(net20),
    .D(_029_),
    .Y(_030_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _117_ (.A(net20),
    .B(_041_),
    .X(_003_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _118_ (.A(net9),
    .B(net8),
    .C(_037_),
    .Y(_031_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _119_ (.A2(_031_),
    .A1(_003_),
    .B1(_030_),
    .X(_001_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _120_ (.A(_030_),
    .B(_031_),
    .X(_002_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _121_ (.Y(_012_),
    .B(_039_),
    .A_N(net46),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _122_ (.A0(net2),
    .A1(net48),
    .S(_039_),
    .X(_013_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _123_ (.Y(_014_),
    .B1(_040_),
    .B2(\mod1.qam16_mod.i_level[3] ),
    .A2(_039_),
    .A1(_035_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dfrbpq_1 _124_ (.RESET_B(net13),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\mod1.qam16_mod.q_level[2] ),
    .Q(\mod1.q_out_qam16[2] ),
    .CLK(clknet_2_0__leaf_clk));
 sg13g2_dfrbpq_1 _125_ (.RESET_B(net13),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\mod1.qam16_mod.q_level[3] ),
    .Q(\mod1.q_out_qam16[3] ),
    .CLK(clknet_2_0__leaf_clk));
 sg13g2_dfrbpq_1 _126_ (.RESET_B(net13),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_009_),
    .Q(\mod1.psk8_mod.q_out[1] ),
    .CLK(clknet_2_2__leaf_clk));
 sg13g2_dfrbpq_1 _127_ (.RESET_B(net13),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_010_),
    .Q(\mod1.psk8_mod.q_out[2] ),
    .CLK(clknet_2_0__leaf_clk));
 sg13g2_dfrbpq_1 _128_ (.RESET_B(net13),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_006_),
    .Q(\mod1.i_out_8psk[0] ),
    .CLK(clknet_2_0__leaf_clk));
 sg13g2_dfrbpq_1 _129_ (.RESET_B(net14),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_007_),
    .Q(\mod1.i_out_8psk[1] ),
    .CLK(clknet_2_3__leaf_clk));
 sg13g2_dfrbpq_1 _130_ (.RESET_B(net15),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_008_),
    .Q(\mod1.i_out_8psk[2] ),
    .CLK(clknet_2_3__leaf_clk));
 sg13g2_dfrbpq_1 _131_ (.RESET_B(net14),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\mod1.qam16_mod.i_level[2] ),
    .Q(\mod1.i_out_qam16[2] ),
    .CLK(clknet_2_1__leaf_clk));
 sg13g2_dfrbpq_1 _132_ (.RESET_B(net15),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\mod1.qam16_mod.i_level[3] ),
    .Q(\mod1.i_out_qam16[3] ),
    .CLK(clknet_2_3__leaf_clk));
 sg13g2_dfrbpq_1 _133_ (.RESET_B(net13),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_012_),
    .Q(\mod1.i_out_qpsk[1] ),
    .CLK(clknet_2_2__leaf_clk));
 sg13g2_dfrbpq_1 _134_ (.RESET_B(net15),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_013_),
    .Q(\mod1.i_out_qpsk[2] ),
    .CLK(clknet_2_2__leaf_clk));
 sg13g2_dfrbpq_1 _135_ (.RESET_B(net14),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_004_),
    .Q(\Demo1.qam16_bits[0] ),
    .CLK(clknet_2_1__leaf_clk));
 sg13g2_dfrbpq_1 _136_ (.RESET_B(net14),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_005_),
    .Q(\Demo1.qam16_bits[1] ),
    .CLK(clknet_2_3__leaf_clk));
 sg13g2_dfrbpq_1 _137_ (.RESET_B(net14),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_011_),
    .Q(\Demo1.qam16_bits[2] ),
    .CLK(clknet_2_1__leaf_clk));
 sg13g2_dfrbpq_1 _138_ (.RESET_B(net14),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_001_),
    .Q(\Demo1.epsk_de1.bit_out[0] ),
    .CLK(clknet_2_1__leaf_clk));
 sg13g2_dfrbpq_1 _139_ (.RESET_B(net15),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_002_),
    .Q(\Demo1.epsk_de1.bit_out[1] ),
    .CLK(clknet_2_3__leaf_clk));
 sg13g2_dfrbpq_1 _140_ (.RESET_B(net14),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_003_),
    .Q(\Demo1.epsk_de1.bit_out[2] ),
    .CLK(clknet_2_1__leaf_clk));
 sg13g2_dfrbpq_1 _141_ (.RESET_B(net13),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_014_),
    .Q(\mod1.q_out_qpsk[2] ),
    .CLK(clknet_2_2__leaf_clk));
 sg13g2_dfrbpq_2 _142_ (.RESET_B(net13),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net37),
    .Q(\Demo1.qam16_bits[3] ),
    .CLK(clknet_2_2__leaf_clk));
 sg13g2_dfrbpq_1 _143_ (.RESET_B(net14),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_000_),
    .Q(\mod1.bpsk_mod.i_out[2] ),
    .CLK(clknet_2_0__leaf_clk));
 sg13g2_tiehi heichips25_template_33 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net38));
 sg13g2_tiehi heichips25_template_34 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net39));
 sg13g2_tiehi heichips25_template_35 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net40));
 sg13g2_tiehi heichips25_template_36 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net41));
 sg13g2_tiehi heichips25_template_37 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net42));
 sg13g2_tiehi heichips25_template_38 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net43));
 sg13g2_tiehi heichips25_template_39 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net44));
 sg13g2_tiehi heichips25_template_40 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net45));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_tielo heichips25_template_29 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net34));
 sg13g2_tielo heichips25_template_30 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net35));
 sg13g2_tielo heichips25_template_31 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net36));
 sg13g2_tiehi _142__32 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net37));
 sg13g2_buf_1 _157_ (.A(net29),
    .X(net25),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout11 (.A(_036_),
    .X(net11),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout12 (.A(_036_),
    .X(net12),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout13 (.A(net15),
    .X(net13),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout14 (.A(net15),
    .X(net14),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout15 (.A(rst_n),
    .X(net15),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 input1 (.A(ui_in[1]),
    .X(net1),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 input2 (.A(ui_in[2]),
    .X(net2),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 input3 (.A(ui_in[3]),
    .X(net3),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 input4 (.A(ui_in[4]),
    .X(net4),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 input5 (.A(ui_in[5]),
    .X(net5),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 input6 (.A(ui_in[6]),
    .X(net6),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 input7 (.A(ui_in[7]),
    .X(net7),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input8 (.A(uio_in[0]),
    .X(net8),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input9 (.A(uio_in[1]),
    .X(net9),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input10 (.A(uio_in[2]),
    .X(net10),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input11 (.A(uio_in[3]),
    .X(net16),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 input12 (.A(uio_in[4]),
    .X(net17),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 input13 (.A(uio_in[5]),
    .X(net18),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 input14 (.A(uio_in[6]),
    .X(net19),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 input15 (.A(uio_in[7]),
    .X(net20),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output16 (.A(net21),
    .X(uio_out[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output17 (.A(net22),
    .X(uio_out[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output18 (.A(net23),
    .X(uio_out[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output19 (.A(net24),
    .X(uio_out[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output20 (.A(net25),
    .X(uo_out[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output21 (.A(net26),
    .X(uo_out[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output22 (.A(net27),
    .X(uo_out[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output23 (.A(net28),
    .X(uo_out[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output24 (.A(net29),
    .X(uo_out[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output25 (.A(net30),
    .X(uo_out[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output26 (.A(net31),
    .X(uo_out[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output27 (.A(net32),
    .X(uo_out[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_tielo heichips25_template_28 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net33));
 sg13g2_buf_8 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 clkload0 (.A(clknet_2_0__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 clkload1 (.A(clknet_2_1__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 clkload2 (.A(clknet_2_3__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlygate4sd3_1 hold1 (.A(\mod1.i_out_qpsk[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net46));
 sg13g2_dlygate4sd3_1 hold2 (.A(\mod1.q_out_qpsk[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net47));
 sg13g2_dlygate4sd3_1 hold3 (.A(\mod1.i_out_qpsk[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net48));
 sg13g2_decap_8 FILLER_0_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_262 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_381 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_479 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_689 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_822 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_370 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_377 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_391 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_412 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_426 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_433 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_440 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_447 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_454 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_475 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_482 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_496 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_503 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_531 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_538 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_615 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_181 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_206 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_213 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_227 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_262 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_381 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_412 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_426 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_433 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_440 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_447 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_454 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_475 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_482 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_496 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_503 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_531 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_538 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_615 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_391 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_446 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_381 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_479 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_689 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_822 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_341 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_348 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_225 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_262 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_381 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_446 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_225 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_232 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_328 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_428 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_435 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_442 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_477 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_596 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_331 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_5 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_12 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_19 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_26 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_33 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_5 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_12 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_19 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_26 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_33 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_414 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_428 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_435 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_442 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_477 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_596 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_5 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_12 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_19 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_26 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_33 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_341 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_348 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_397 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_446 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_5 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_12 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_19 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_26 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_33 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_446 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_5 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_12 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_19 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_26 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_33 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_331 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_391 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_412 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_426 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_433 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_440 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_447 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_454 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_475 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_482 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_496 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_503 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_531 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_538 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_615 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_5 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_12 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_19 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_26 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_33 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_262 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_381 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_479 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_689 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_822 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_5 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_12 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_19 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_26 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_33 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_328 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_370 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_377 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_391 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_412 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_426 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_433 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_440 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_447 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_454 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_475 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_482 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_496 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_503 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_531 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_538 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_615 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_414 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_428 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_435 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_442 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_477 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_596 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_341 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_348 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_397 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_446 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_341 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_348 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_397 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_446 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_5 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_12 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_19 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_26 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_33 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_341 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_348 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_397 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_446 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_5 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_12 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_19 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_26 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_33 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_341 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_348 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_397 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_446 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_5 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_12 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_19 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_26 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_33 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_341 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_348 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_397 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_446 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_5 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_12 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_19 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_26 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_33 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_341 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_348 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_397 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_446 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_1022 (.VDD(VPWR),
    .VSS(VGND));
 assign uio_oe[0] = net38;
 assign uio_oe[1] = net39;
 assign uio_oe[2] = net40;
 assign uio_oe[3] = net41;
 assign uio_oe[4] = net42;
 assign uio_oe[5] = net43;
 assign uio_oe[6] = net44;
 assign uio_oe[7] = net45;
 assign uio_out[4] = net33;
 assign uio_out[5] = net34;
 assign uio_out[6] = net35;
 assign uio_out[7] = net36;
endmodule
