magic
tech ihp-sg13g2
magscale 1 2
timestamp 1754656326
<< metal1 >>
rect 576 38576 99360 38600
rect 576 38536 4352 38576
rect 4392 38536 4434 38576
rect 4474 38536 4516 38576
rect 4556 38536 4598 38576
rect 4638 38536 4680 38576
rect 4720 38536 19472 38576
rect 19512 38536 19554 38576
rect 19594 38536 19636 38576
rect 19676 38536 19718 38576
rect 19758 38536 19800 38576
rect 19840 38536 34592 38576
rect 34632 38536 34674 38576
rect 34714 38536 34756 38576
rect 34796 38536 34838 38576
rect 34878 38536 34920 38576
rect 34960 38536 49712 38576
rect 49752 38536 49794 38576
rect 49834 38536 49876 38576
rect 49916 38536 49958 38576
rect 49998 38536 50040 38576
rect 50080 38536 64832 38576
rect 64872 38536 64914 38576
rect 64954 38536 64996 38576
rect 65036 38536 65078 38576
rect 65118 38536 65160 38576
rect 65200 38536 79952 38576
rect 79992 38536 80034 38576
rect 80074 38536 80116 38576
rect 80156 38536 80198 38576
rect 80238 38536 80280 38576
rect 80320 38536 95072 38576
rect 95112 38536 95154 38576
rect 95194 38536 95236 38576
rect 95276 38536 95318 38576
rect 95358 38536 95400 38576
rect 95440 38536 99360 38576
rect 576 38512 99360 38536
rect 576 37820 99360 37844
rect 576 37780 3112 37820
rect 3152 37780 3194 37820
rect 3234 37780 3276 37820
rect 3316 37780 3358 37820
rect 3398 37780 3440 37820
rect 3480 37780 18232 37820
rect 18272 37780 18314 37820
rect 18354 37780 18396 37820
rect 18436 37780 18478 37820
rect 18518 37780 18560 37820
rect 18600 37780 33352 37820
rect 33392 37780 33434 37820
rect 33474 37780 33516 37820
rect 33556 37780 33598 37820
rect 33638 37780 33680 37820
rect 33720 37780 48472 37820
rect 48512 37780 48554 37820
rect 48594 37780 48636 37820
rect 48676 37780 48718 37820
rect 48758 37780 48800 37820
rect 48840 37780 63592 37820
rect 63632 37780 63674 37820
rect 63714 37780 63756 37820
rect 63796 37780 63838 37820
rect 63878 37780 63920 37820
rect 63960 37780 78712 37820
rect 78752 37780 78794 37820
rect 78834 37780 78876 37820
rect 78916 37780 78958 37820
rect 78998 37780 79040 37820
rect 79080 37780 93832 37820
rect 93872 37780 93914 37820
rect 93954 37780 93996 37820
rect 94036 37780 94078 37820
rect 94118 37780 94160 37820
rect 94200 37780 99360 37820
rect 576 37756 99360 37780
rect 576 37064 99360 37088
rect 576 37024 4352 37064
rect 4392 37024 4434 37064
rect 4474 37024 4516 37064
rect 4556 37024 4598 37064
rect 4638 37024 4680 37064
rect 4720 37024 19472 37064
rect 19512 37024 19554 37064
rect 19594 37024 19636 37064
rect 19676 37024 19718 37064
rect 19758 37024 19800 37064
rect 19840 37024 34592 37064
rect 34632 37024 34674 37064
rect 34714 37024 34756 37064
rect 34796 37024 34838 37064
rect 34878 37024 34920 37064
rect 34960 37024 49712 37064
rect 49752 37024 49794 37064
rect 49834 37024 49876 37064
rect 49916 37024 49958 37064
rect 49998 37024 50040 37064
rect 50080 37024 64832 37064
rect 64872 37024 64914 37064
rect 64954 37024 64996 37064
rect 65036 37024 65078 37064
rect 65118 37024 65160 37064
rect 65200 37024 79952 37064
rect 79992 37024 80034 37064
rect 80074 37024 80116 37064
rect 80156 37024 80198 37064
rect 80238 37024 80280 37064
rect 80320 37024 95072 37064
rect 95112 37024 95154 37064
rect 95194 37024 95236 37064
rect 95276 37024 95318 37064
rect 95358 37024 95400 37064
rect 95440 37024 99360 37064
rect 576 37000 99360 37024
rect 576 36308 99360 36332
rect 576 36268 3112 36308
rect 3152 36268 3194 36308
rect 3234 36268 3276 36308
rect 3316 36268 3358 36308
rect 3398 36268 3440 36308
rect 3480 36268 18232 36308
rect 18272 36268 18314 36308
rect 18354 36268 18396 36308
rect 18436 36268 18478 36308
rect 18518 36268 18560 36308
rect 18600 36268 33352 36308
rect 33392 36268 33434 36308
rect 33474 36268 33516 36308
rect 33556 36268 33598 36308
rect 33638 36268 33680 36308
rect 33720 36268 48472 36308
rect 48512 36268 48554 36308
rect 48594 36268 48636 36308
rect 48676 36268 48718 36308
rect 48758 36268 48800 36308
rect 48840 36268 63592 36308
rect 63632 36268 63674 36308
rect 63714 36268 63756 36308
rect 63796 36268 63838 36308
rect 63878 36268 63920 36308
rect 63960 36268 78712 36308
rect 78752 36268 78794 36308
rect 78834 36268 78876 36308
rect 78916 36268 78958 36308
rect 78998 36268 79040 36308
rect 79080 36268 93832 36308
rect 93872 36268 93914 36308
rect 93954 36268 93996 36308
rect 94036 36268 94078 36308
rect 94118 36268 94160 36308
rect 94200 36268 99360 36308
rect 576 36244 99360 36268
rect 576 35552 99360 35576
rect 576 35512 4352 35552
rect 4392 35512 4434 35552
rect 4474 35512 4516 35552
rect 4556 35512 4598 35552
rect 4638 35512 4680 35552
rect 4720 35512 19472 35552
rect 19512 35512 19554 35552
rect 19594 35512 19636 35552
rect 19676 35512 19718 35552
rect 19758 35512 19800 35552
rect 19840 35512 34592 35552
rect 34632 35512 34674 35552
rect 34714 35512 34756 35552
rect 34796 35512 34838 35552
rect 34878 35512 34920 35552
rect 34960 35512 49712 35552
rect 49752 35512 49794 35552
rect 49834 35512 49876 35552
rect 49916 35512 49958 35552
rect 49998 35512 50040 35552
rect 50080 35512 64832 35552
rect 64872 35512 64914 35552
rect 64954 35512 64996 35552
rect 65036 35512 65078 35552
rect 65118 35512 65160 35552
rect 65200 35512 79952 35552
rect 79992 35512 80034 35552
rect 80074 35512 80116 35552
rect 80156 35512 80198 35552
rect 80238 35512 80280 35552
rect 80320 35512 95072 35552
rect 95112 35512 95154 35552
rect 95194 35512 95236 35552
rect 95276 35512 95318 35552
rect 95358 35512 95400 35552
rect 95440 35512 99360 35552
rect 576 35488 99360 35512
rect 643 35216 701 35217
rect 643 35176 652 35216
rect 692 35176 701 35216
rect 643 35175 701 35176
rect 835 35216 893 35217
rect 835 35176 844 35216
rect 884 35176 893 35216
rect 835 35175 893 35176
rect 576 34796 99360 34820
rect 576 34756 3112 34796
rect 3152 34756 3194 34796
rect 3234 34756 3276 34796
rect 3316 34756 3358 34796
rect 3398 34756 3440 34796
rect 3480 34756 18232 34796
rect 18272 34756 18314 34796
rect 18354 34756 18396 34796
rect 18436 34756 18478 34796
rect 18518 34756 18560 34796
rect 18600 34756 33352 34796
rect 33392 34756 33434 34796
rect 33474 34756 33516 34796
rect 33556 34756 33598 34796
rect 33638 34756 33680 34796
rect 33720 34756 48472 34796
rect 48512 34756 48554 34796
rect 48594 34756 48636 34796
rect 48676 34756 48718 34796
rect 48758 34756 48800 34796
rect 48840 34756 63592 34796
rect 63632 34756 63674 34796
rect 63714 34756 63756 34796
rect 63796 34756 63838 34796
rect 63878 34756 63920 34796
rect 63960 34756 78712 34796
rect 78752 34756 78794 34796
rect 78834 34756 78876 34796
rect 78916 34756 78958 34796
rect 78998 34756 79040 34796
rect 79080 34756 93832 34796
rect 93872 34756 93914 34796
rect 93954 34756 93996 34796
rect 94036 34756 94078 34796
rect 94118 34756 94160 34796
rect 94200 34756 99360 34796
rect 576 34732 99360 34756
rect 643 34376 701 34377
rect 643 34336 652 34376
rect 692 34336 701 34376
rect 643 34335 701 34336
rect 835 34376 893 34377
rect 835 34336 844 34376
rect 884 34336 893 34376
rect 835 34335 893 34336
rect 576 34040 99360 34064
rect 576 34000 4352 34040
rect 4392 34000 4434 34040
rect 4474 34000 4516 34040
rect 4556 34000 4598 34040
rect 4638 34000 4680 34040
rect 4720 34000 19472 34040
rect 19512 34000 19554 34040
rect 19594 34000 19636 34040
rect 19676 34000 19718 34040
rect 19758 34000 19800 34040
rect 19840 34000 34592 34040
rect 34632 34000 34674 34040
rect 34714 34000 34756 34040
rect 34796 34000 34838 34040
rect 34878 34000 34920 34040
rect 34960 34000 49712 34040
rect 49752 34000 49794 34040
rect 49834 34000 49876 34040
rect 49916 34000 49958 34040
rect 49998 34000 50040 34040
rect 50080 34000 64832 34040
rect 64872 34000 64914 34040
rect 64954 34000 64996 34040
rect 65036 34000 65078 34040
rect 65118 34000 65160 34040
rect 65200 34000 79952 34040
rect 79992 34000 80034 34040
rect 80074 34000 80116 34040
rect 80156 34000 80198 34040
rect 80238 34000 80280 34040
rect 80320 34000 95072 34040
rect 95112 34000 95154 34040
rect 95194 34000 95236 34040
rect 95276 34000 95318 34040
rect 95358 34000 95400 34040
rect 95440 34000 99360 34040
rect 576 33976 99360 34000
rect 643 33704 701 33705
rect 643 33664 652 33704
rect 692 33664 701 33704
rect 643 33663 701 33664
rect 835 33704 893 33705
rect 835 33664 844 33704
rect 884 33664 893 33704
rect 835 33663 893 33664
rect 576 33284 99360 33308
rect 576 33244 3112 33284
rect 3152 33244 3194 33284
rect 3234 33244 3276 33284
rect 3316 33244 3358 33284
rect 3398 33244 3440 33284
rect 3480 33244 18232 33284
rect 18272 33244 18314 33284
rect 18354 33244 18396 33284
rect 18436 33244 18478 33284
rect 18518 33244 18560 33284
rect 18600 33244 33352 33284
rect 33392 33244 33434 33284
rect 33474 33244 33516 33284
rect 33556 33244 33598 33284
rect 33638 33244 33680 33284
rect 33720 33244 48472 33284
rect 48512 33244 48554 33284
rect 48594 33244 48636 33284
rect 48676 33244 48718 33284
rect 48758 33244 48800 33284
rect 48840 33244 63592 33284
rect 63632 33244 63674 33284
rect 63714 33244 63756 33284
rect 63796 33244 63838 33284
rect 63878 33244 63920 33284
rect 63960 33244 78712 33284
rect 78752 33244 78794 33284
rect 78834 33244 78876 33284
rect 78916 33244 78958 33284
rect 78998 33244 79040 33284
rect 79080 33244 93832 33284
rect 93872 33244 93914 33284
rect 93954 33244 93996 33284
rect 94036 33244 94078 33284
rect 94118 33244 94160 33284
rect 94200 33244 99360 33284
rect 576 33220 99360 33244
rect 643 32864 701 32865
rect 643 32824 652 32864
rect 692 32824 701 32864
rect 643 32823 701 32824
rect 835 32864 893 32865
rect 835 32824 844 32864
rect 884 32824 893 32864
rect 835 32823 893 32824
rect 576 32528 99360 32552
rect 576 32488 4352 32528
rect 4392 32488 4434 32528
rect 4474 32488 4516 32528
rect 4556 32488 4598 32528
rect 4638 32488 4680 32528
rect 4720 32488 19472 32528
rect 19512 32488 19554 32528
rect 19594 32488 19636 32528
rect 19676 32488 19718 32528
rect 19758 32488 19800 32528
rect 19840 32488 34592 32528
rect 34632 32488 34674 32528
rect 34714 32488 34756 32528
rect 34796 32488 34838 32528
rect 34878 32488 34920 32528
rect 34960 32488 49712 32528
rect 49752 32488 49794 32528
rect 49834 32488 49876 32528
rect 49916 32488 49958 32528
rect 49998 32488 50040 32528
rect 50080 32488 64832 32528
rect 64872 32488 64914 32528
rect 64954 32488 64996 32528
rect 65036 32488 65078 32528
rect 65118 32488 65160 32528
rect 65200 32488 79952 32528
rect 79992 32488 80034 32528
rect 80074 32488 80116 32528
rect 80156 32488 80198 32528
rect 80238 32488 80280 32528
rect 80320 32488 95072 32528
rect 95112 32488 95154 32528
rect 95194 32488 95236 32528
rect 95276 32488 95318 32528
rect 95358 32488 95400 32528
rect 95440 32488 99360 32528
rect 576 32464 99360 32488
rect 27435 32192 27477 32201
rect 27435 32152 27436 32192
rect 27476 32152 27477 32192
rect 27435 32143 27477 32152
rect 643 32108 701 32109
rect 643 32068 652 32108
rect 692 32068 701 32108
rect 643 32067 701 32068
rect 843 31940 885 31949
rect 843 31900 844 31940
rect 884 31900 885 31940
rect 843 31891 885 31900
rect 27531 31940 27573 31949
rect 27531 31900 27532 31940
rect 27572 31900 27573 31940
rect 27531 31891 27573 31900
rect 576 31772 99360 31796
rect 576 31732 3112 31772
rect 3152 31732 3194 31772
rect 3234 31732 3276 31772
rect 3316 31732 3358 31772
rect 3398 31732 3440 31772
rect 3480 31732 18232 31772
rect 18272 31732 18314 31772
rect 18354 31732 18396 31772
rect 18436 31732 18478 31772
rect 18518 31732 18560 31772
rect 18600 31732 33352 31772
rect 33392 31732 33434 31772
rect 33474 31732 33516 31772
rect 33556 31732 33598 31772
rect 33638 31732 33680 31772
rect 33720 31732 48472 31772
rect 48512 31732 48554 31772
rect 48594 31732 48636 31772
rect 48676 31732 48718 31772
rect 48758 31732 48800 31772
rect 48840 31732 63592 31772
rect 63632 31732 63674 31772
rect 63714 31732 63756 31772
rect 63796 31732 63838 31772
rect 63878 31732 63920 31772
rect 63960 31732 78712 31772
rect 78752 31732 78794 31772
rect 78834 31732 78876 31772
rect 78916 31732 78958 31772
rect 78998 31732 79040 31772
rect 79080 31732 93832 31772
rect 93872 31732 93914 31772
rect 93954 31732 93996 31772
rect 94036 31732 94078 31772
rect 94118 31732 94160 31772
rect 94200 31732 99360 31772
rect 576 31708 99360 31732
rect 643 31436 701 31437
rect 643 31396 652 31436
rect 692 31396 701 31436
rect 643 31395 701 31396
rect 21763 31352 21821 31353
rect 21763 31312 21772 31352
rect 21812 31312 21821 31352
rect 21763 31311 21821 31312
rect 22627 31352 22685 31353
rect 22627 31312 22636 31352
rect 22676 31312 22685 31352
rect 22627 31311 22685 31312
rect 27907 31352 27965 31353
rect 27907 31312 27916 31352
rect 27956 31312 27965 31352
rect 27907 31311 27965 31312
rect 28771 31352 28829 31353
rect 28771 31312 28780 31352
rect 28820 31312 28829 31352
rect 28771 31311 28829 31312
rect 21387 31268 21429 31277
rect 21387 31228 21388 31268
rect 21428 31228 21429 31268
rect 21387 31219 21429 31228
rect 29163 31268 29205 31277
rect 29163 31228 29164 31268
rect 29204 31228 29205 31268
rect 29163 31219 29205 31228
rect 843 31184 885 31193
rect 843 31144 844 31184
rect 884 31144 885 31184
rect 843 31135 885 31144
rect 23779 31184 23837 31185
rect 23779 31144 23788 31184
rect 23828 31144 23837 31184
rect 23779 31143 23837 31144
rect 26755 31184 26813 31185
rect 26755 31144 26764 31184
rect 26804 31144 26813 31184
rect 26755 31143 26813 31144
rect 576 31016 99360 31040
rect 576 30976 4352 31016
rect 4392 30976 4434 31016
rect 4474 30976 4516 31016
rect 4556 30976 4598 31016
rect 4638 30976 4680 31016
rect 4720 30976 19472 31016
rect 19512 30976 19554 31016
rect 19594 30976 19636 31016
rect 19676 30976 19718 31016
rect 19758 30976 19800 31016
rect 19840 30976 34592 31016
rect 34632 30976 34674 31016
rect 34714 30976 34756 31016
rect 34796 30976 34838 31016
rect 34878 30976 34920 31016
rect 34960 30976 49712 31016
rect 49752 30976 49794 31016
rect 49834 30976 49876 31016
rect 49916 30976 49958 31016
rect 49998 30976 50040 31016
rect 50080 30976 64832 31016
rect 64872 30976 64914 31016
rect 64954 30976 64996 31016
rect 65036 30976 65078 31016
rect 65118 30976 65160 31016
rect 65200 30976 79952 31016
rect 79992 30976 80034 31016
rect 80074 30976 80116 31016
rect 80156 30976 80198 31016
rect 80238 30976 80280 31016
rect 80320 30976 95072 31016
rect 95112 30976 95154 31016
rect 95194 30976 95236 31016
rect 95276 30976 95318 31016
rect 95358 30976 95400 31016
rect 95440 30976 99360 31016
rect 576 30952 99360 30976
rect 27243 30680 27285 30689
rect 27243 30640 27244 30680
rect 27284 30640 27285 30680
rect 27243 30631 27285 30640
rect 27619 30680 27677 30681
rect 27619 30640 27628 30680
rect 27668 30640 27677 30680
rect 27619 30639 27677 30640
rect 32715 30680 32757 30689
rect 32715 30640 32716 30680
rect 32756 30640 32757 30680
rect 32715 30631 32757 30640
rect 33091 30680 33149 30681
rect 33091 30640 33100 30680
rect 33140 30640 33149 30680
rect 33091 30639 33149 30640
rect 33955 30680 34013 30681
rect 33955 30640 33964 30680
rect 34004 30640 34013 30680
rect 33955 30639 34013 30640
rect 643 30596 701 30597
rect 643 30556 652 30596
rect 692 30556 701 30596
rect 643 30555 701 30556
rect 27339 30596 27381 30605
rect 27339 30556 27340 30596
rect 27380 30556 27381 30596
rect 27339 30547 27381 30556
rect 27531 30596 27573 30605
rect 27531 30556 27532 30596
rect 27572 30556 27573 30596
rect 27531 30547 27573 30556
rect 27435 30512 27477 30521
rect 27435 30472 27436 30512
rect 27476 30472 27477 30512
rect 27435 30463 27477 30472
rect 843 30428 885 30437
rect 843 30388 844 30428
rect 884 30388 885 30428
rect 843 30379 885 30388
rect 35107 30428 35165 30429
rect 35107 30388 35116 30428
rect 35156 30388 35165 30428
rect 35107 30387 35165 30388
rect 576 30260 99360 30284
rect 576 30220 3112 30260
rect 3152 30220 3194 30260
rect 3234 30220 3276 30260
rect 3316 30220 3358 30260
rect 3398 30220 3440 30260
rect 3480 30220 18232 30260
rect 18272 30220 18314 30260
rect 18354 30220 18396 30260
rect 18436 30220 18478 30260
rect 18518 30220 18560 30260
rect 18600 30220 33352 30260
rect 33392 30220 33434 30260
rect 33474 30220 33516 30260
rect 33556 30220 33598 30260
rect 33638 30220 33680 30260
rect 33720 30220 48472 30260
rect 48512 30220 48554 30260
rect 48594 30220 48636 30260
rect 48676 30220 48718 30260
rect 48758 30220 48800 30260
rect 48840 30220 63592 30260
rect 63632 30220 63674 30260
rect 63714 30220 63756 30260
rect 63796 30220 63838 30260
rect 63878 30220 63920 30260
rect 63960 30220 78712 30260
rect 78752 30220 78794 30260
rect 78834 30220 78876 30260
rect 78916 30220 78958 30260
rect 78998 30220 79040 30260
rect 79080 30220 93832 30260
rect 93872 30220 93914 30260
rect 93954 30220 93996 30260
rect 94036 30220 94078 30260
rect 94118 30220 94160 30260
rect 94200 30220 99360 30260
rect 576 30196 99360 30220
rect 643 29924 701 29925
rect 643 29884 652 29924
rect 692 29884 701 29924
rect 643 29883 701 29884
rect 36459 29840 36501 29849
rect 36459 29800 36460 29840
rect 36500 29800 36501 29840
rect 36459 29791 36501 29800
rect 843 29672 885 29681
rect 843 29632 844 29672
rect 884 29632 885 29672
rect 843 29623 885 29632
rect 36747 29672 36789 29681
rect 36747 29632 36748 29672
rect 36788 29632 36789 29672
rect 36747 29623 36789 29632
rect 576 29504 99360 29528
rect 576 29464 4352 29504
rect 4392 29464 4434 29504
rect 4474 29464 4516 29504
rect 4556 29464 4598 29504
rect 4638 29464 4680 29504
rect 4720 29464 19472 29504
rect 19512 29464 19554 29504
rect 19594 29464 19636 29504
rect 19676 29464 19718 29504
rect 19758 29464 19800 29504
rect 19840 29464 34592 29504
rect 34632 29464 34674 29504
rect 34714 29464 34756 29504
rect 34796 29464 34838 29504
rect 34878 29464 34920 29504
rect 34960 29464 49712 29504
rect 49752 29464 49794 29504
rect 49834 29464 49876 29504
rect 49916 29464 49958 29504
rect 49998 29464 50040 29504
rect 50080 29464 64832 29504
rect 64872 29464 64914 29504
rect 64954 29464 64996 29504
rect 65036 29464 65078 29504
rect 65118 29464 65160 29504
rect 65200 29464 79952 29504
rect 79992 29464 80034 29504
rect 80074 29464 80116 29504
rect 80156 29464 80198 29504
rect 80238 29464 80280 29504
rect 80320 29464 95072 29504
rect 95112 29464 95154 29504
rect 95194 29464 95236 29504
rect 95276 29464 95318 29504
rect 95358 29464 95400 29504
rect 95440 29464 99360 29504
rect 576 29440 99360 29464
rect 31275 29336 31317 29345
rect 31275 29296 31276 29336
rect 31316 29296 31317 29336
rect 31275 29287 31317 29296
rect 15339 29168 15381 29177
rect 15339 29128 15340 29168
rect 15380 29128 15381 29168
rect 15339 29119 15381 29128
rect 15715 29168 15773 29169
rect 15715 29128 15724 29168
rect 15764 29128 15773 29168
rect 15715 29127 15773 29128
rect 16579 29168 16637 29169
rect 16579 29128 16588 29168
rect 16628 29128 16637 29168
rect 16579 29127 16637 29128
rect 31171 29168 31229 29169
rect 31171 29128 31180 29168
rect 31220 29128 31229 29168
rect 31171 29127 31229 29128
rect 35587 29168 35645 29169
rect 35587 29128 35596 29168
rect 35636 29128 35645 29168
rect 35587 29127 35645 29128
rect 35979 29168 36021 29177
rect 35979 29128 35980 29168
rect 36020 29128 36021 29168
rect 35979 29119 36021 29128
rect 35691 29084 35733 29093
rect 35691 29044 35692 29084
rect 35732 29044 35733 29084
rect 35691 29035 35733 29044
rect 35883 29084 35925 29093
rect 35883 29044 35884 29084
rect 35924 29044 35925 29084
rect 35883 29035 35925 29044
rect 35787 29000 35829 29009
rect 35787 28960 35788 29000
rect 35828 28960 35829 29000
rect 35787 28951 35829 28960
rect 17731 28916 17789 28917
rect 17731 28876 17740 28916
rect 17780 28876 17789 28916
rect 17731 28875 17789 28876
rect 576 28748 99360 28772
rect 576 28708 3112 28748
rect 3152 28708 3194 28748
rect 3234 28708 3276 28748
rect 3316 28708 3358 28748
rect 3398 28708 3440 28748
rect 3480 28708 18232 28748
rect 18272 28708 18314 28748
rect 18354 28708 18396 28748
rect 18436 28708 18478 28748
rect 18518 28708 18560 28748
rect 18600 28708 33352 28748
rect 33392 28708 33434 28748
rect 33474 28708 33516 28748
rect 33556 28708 33598 28748
rect 33638 28708 33680 28748
rect 33720 28708 48472 28748
rect 48512 28708 48554 28748
rect 48594 28708 48636 28748
rect 48676 28708 48718 28748
rect 48758 28708 48800 28748
rect 48840 28708 63592 28748
rect 63632 28708 63674 28748
rect 63714 28708 63756 28748
rect 63796 28708 63838 28748
rect 63878 28708 63920 28748
rect 63960 28708 78712 28748
rect 78752 28708 78794 28748
rect 78834 28708 78876 28748
rect 78916 28708 78958 28748
rect 78998 28708 79040 28748
rect 79080 28708 93832 28748
rect 93872 28708 93914 28748
rect 93954 28708 93996 28748
rect 94036 28708 94078 28748
rect 94118 28708 94160 28748
rect 94200 28708 99360 28748
rect 576 28684 99360 28708
rect 22059 28580 22101 28589
rect 22059 28540 22060 28580
rect 22100 28540 22101 28580
rect 22059 28531 22101 28540
rect 28299 28496 28341 28505
rect 28299 28456 28300 28496
rect 28340 28456 28341 28496
rect 28299 28447 28341 28456
rect 28779 28496 28821 28505
rect 28779 28456 28780 28496
rect 28820 28456 28821 28496
rect 28779 28447 28821 28456
rect 28203 28412 28245 28421
rect 28203 28372 28204 28412
rect 28244 28372 28245 28412
rect 28203 28363 28245 28372
rect 28395 28412 28437 28421
rect 28395 28372 28396 28412
rect 28436 28372 28437 28412
rect 28395 28363 28437 28372
rect 643 28328 701 28329
rect 643 28288 652 28328
rect 692 28288 701 28328
rect 643 28287 701 28288
rect 835 28328 893 28329
rect 835 28288 844 28328
rect 884 28288 893 28328
rect 835 28287 893 28288
rect 22347 28328 22389 28337
rect 22347 28288 22348 28328
rect 22388 28288 22389 28328
rect 22347 28279 22389 28288
rect 22435 28328 22493 28329
rect 22435 28288 22444 28328
rect 22484 28288 22493 28328
rect 22435 28287 22493 28288
rect 23395 28328 23453 28329
rect 23395 28288 23404 28328
rect 23444 28288 23453 28328
rect 23395 28287 23453 28288
rect 28099 28328 28157 28329
rect 28099 28288 28108 28328
rect 28148 28288 28157 28328
rect 28099 28287 28157 28288
rect 28491 28328 28533 28337
rect 28491 28288 28492 28328
rect 28532 28288 28533 28328
rect 28491 28279 28533 28288
rect 29067 28328 29109 28337
rect 29067 28288 29068 28328
rect 29108 28288 29109 28328
rect 29067 28279 29109 28288
rect 29155 28328 29213 28329
rect 29155 28288 29164 28328
rect 29204 28288 29213 28328
rect 29155 28287 29213 28288
rect 29443 28328 29501 28329
rect 29443 28288 29452 28328
rect 29492 28288 29501 28328
rect 29443 28287 29501 28288
rect 29643 28328 29685 28337
rect 29643 28288 29644 28328
rect 29684 28288 29685 28328
rect 29643 28279 29685 28288
rect 29731 28328 29789 28329
rect 29731 28288 29740 28328
rect 29780 28288 29789 28328
rect 29731 28287 29789 28288
rect 23203 28244 23261 28245
rect 23203 28204 23212 28244
rect 23252 28204 23261 28244
rect 23203 28203 23261 28204
rect 23491 28160 23549 28161
rect 23491 28120 23500 28160
rect 23540 28120 23549 28160
rect 23491 28119 23549 28120
rect 29451 28160 29493 28169
rect 29451 28120 29452 28160
rect 29492 28120 29493 28160
rect 29451 28111 29493 28120
rect 22539 28102 22581 28111
rect 22539 28062 22540 28102
rect 22580 28062 22581 28102
rect 22539 28053 22581 28062
rect 29259 28102 29301 28111
rect 29259 28062 29260 28102
rect 29300 28062 29301 28102
rect 29259 28053 29301 28062
rect 576 27992 99360 28016
rect 576 27952 4352 27992
rect 4392 27952 4434 27992
rect 4474 27952 4516 27992
rect 4556 27952 4598 27992
rect 4638 27952 4680 27992
rect 4720 27952 19472 27992
rect 19512 27952 19554 27992
rect 19594 27952 19636 27992
rect 19676 27952 19718 27992
rect 19758 27952 19800 27992
rect 19840 27952 34592 27992
rect 34632 27952 34674 27992
rect 34714 27952 34756 27992
rect 34796 27952 34838 27992
rect 34878 27952 34920 27992
rect 34960 27952 49712 27992
rect 49752 27952 49794 27992
rect 49834 27952 49876 27992
rect 49916 27952 49958 27992
rect 49998 27952 50040 27992
rect 50080 27952 64832 27992
rect 64872 27952 64914 27992
rect 64954 27952 64996 27992
rect 65036 27952 65078 27992
rect 65118 27952 65160 27992
rect 65200 27952 79952 27992
rect 79992 27952 80034 27992
rect 80074 27952 80116 27992
rect 80156 27952 80198 27992
rect 80238 27952 80280 27992
rect 80320 27952 95072 27992
rect 95112 27952 95154 27992
rect 95194 27952 95236 27992
rect 95276 27952 95318 27992
rect 95358 27952 95400 27992
rect 95440 27952 99360 27992
rect 576 27928 99360 27952
rect 20035 27824 20093 27825
rect 20035 27784 20044 27824
rect 20084 27784 20093 27824
rect 20035 27783 20093 27784
rect 23299 27824 23357 27825
rect 23299 27784 23308 27824
rect 23348 27784 23357 27824
rect 23299 27783 23357 27784
rect 26851 27824 26909 27825
rect 26851 27784 26860 27824
rect 26900 27784 26909 27824
rect 26851 27783 26909 27784
rect 26571 27740 26613 27749
rect 26571 27700 26572 27740
rect 26612 27700 26613 27740
rect 26571 27691 26613 27700
rect 27139 27740 27197 27741
rect 27139 27700 27148 27740
rect 27188 27700 27197 27740
rect 27139 27699 27197 27700
rect 643 27656 701 27657
rect 643 27616 652 27656
rect 692 27616 701 27656
rect 643 27615 701 27616
rect 835 27656 893 27657
rect 835 27616 844 27656
rect 884 27616 893 27656
rect 835 27615 893 27616
rect 18115 27656 18173 27657
rect 18115 27616 18124 27656
rect 18164 27616 18173 27656
rect 18115 27615 18173 27616
rect 18507 27656 18549 27665
rect 18507 27616 18508 27656
rect 18548 27616 18549 27656
rect 18507 27607 18549 27616
rect 18691 27656 18749 27657
rect 18691 27616 18700 27656
rect 18740 27616 18749 27656
rect 18691 27615 18749 27616
rect 20131 27656 20189 27657
rect 20131 27616 20140 27656
rect 20180 27616 20189 27656
rect 20131 27615 20189 27616
rect 23395 27656 23453 27657
rect 23395 27616 23404 27656
rect 23444 27616 23453 27656
rect 23395 27615 23453 27616
rect 26379 27656 26421 27665
rect 26379 27616 26380 27656
rect 26420 27616 26421 27656
rect 26379 27607 26421 27616
rect 26667 27656 26709 27665
rect 26667 27616 26668 27656
rect 26708 27616 26709 27656
rect 26667 27607 26709 27616
rect 26947 27656 27005 27657
rect 26947 27616 26956 27656
rect 26996 27616 27005 27656
rect 26947 27615 27005 27616
rect 29547 27656 29589 27665
rect 29547 27616 29548 27656
rect 29588 27616 29589 27656
rect 29547 27607 29589 27616
rect 29635 27640 29693 27641
rect 29635 27600 29644 27640
rect 29684 27600 29693 27640
rect 29635 27599 29693 27600
rect 18219 27572 18261 27581
rect 18219 27532 18220 27572
rect 18260 27532 18261 27572
rect 18219 27523 18261 27532
rect 18411 27572 18453 27581
rect 18411 27532 18412 27572
rect 18452 27532 18453 27572
rect 18411 27523 18453 27532
rect 29451 27572 29493 27581
rect 29451 27532 29452 27572
rect 29492 27532 29493 27572
rect 29451 27523 29493 27532
rect 18315 27488 18357 27497
rect 18315 27448 18316 27488
rect 18356 27448 18357 27488
rect 18315 27439 18357 27448
rect 29259 27488 29301 27497
rect 29259 27448 29260 27488
rect 29300 27448 29301 27488
rect 29259 27439 29301 27448
rect 29347 27446 29405 27447
rect 18795 27404 18837 27413
rect 29347 27406 29356 27446
rect 29396 27406 29405 27446
rect 29347 27405 29405 27406
rect 18795 27364 18796 27404
rect 18836 27364 18837 27404
rect 18795 27355 18837 27364
rect 20323 27404 20381 27405
rect 20323 27364 20332 27404
rect 20372 27364 20381 27404
rect 20323 27363 20381 27364
rect 23587 27404 23645 27405
rect 23587 27364 23596 27404
rect 23636 27364 23645 27404
rect 23587 27363 23645 27364
rect 576 27236 99360 27260
rect 576 27196 3112 27236
rect 3152 27196 3194 27236
rect 3234 27196 3276 27236
rect 3316 27196 3358 27236
rect 3398 27196 3440 27236
rect 3480 27196 18232 27236
rect 18272 27196 18314 27236
rect 18354 27196 18396 27236
rect 18436 27196 18478 27236
rect 18518 27196 18560 27236
rect 18600 27196 33352 27236
rect 33392 27196 33434 27236
rect 33474 27196 33516 27236
rect 33556 27196 33598 27236
rect 33638 27196 33680 27236
rect 33720 27196 48472 27236
rect 48512 27196 48554 27236
rect 48594 27196 48636 27236
rect 48676 27196 48718 27236
rect 48758 27196 48800 27236
rect 48840 27196 63592 27236
rect 63632 27196 63674 27236
rect 63714 27196 63756 27236
rect 63796 27196 63838 27236
rect 63878 27196 63920 27236
rect 63960 27196 78712 27236
rect 78752 27196 78794 27236
rect 78834 27196 78876 27236
rect 78916 27196 78958 27236
rect 78998 27196 79040 27236
rect 79080 27196 93832 27236
rect 93872 27196 93914 27236
rect 93954 27196 93996 27236
rect 94036 27196 94078 27236
rect 94118 27196 94160 27236
rect 94200 27196 99360 27236
rect 576 27172 99360 27196
rect 29451 27068 29493 27077
rect 29451 27028 29452 27068
rect 29492 27028 29493 27068
rect 29451 27019 29493 27028
rect 29931 27068 29973 27077
rect 29931 27028 29932 27068
rect 29972 27028 29973 27068
rect 29931 27019 29973 27028
rect 37315 27068 37373 27069
rect 37315 27028 37324 27068
rect 37364 27028 37373 27068
rect 37315 27027 37373 27028
rect 19947 26984 19989 26993
rect 19947 26944 19948 26984
rect 19988 26944 19989 26984
rect 19947 26935 19989 26944
rect 29643 26984 29685 26993
rect 29643 26944 29644 26984
rect 29684 26944 29685 26984
rect 29643 26935 29685 26944
rect 30123 26984 30165 26993
rect 30123 26944 30124 26984
rect 30164 26944 30165 26984
rect 30123 26935 30165 26944
rect 643 26816 701 26817
rect 643 26776 652 26816
rect 692 26776 701 26816
rect 643 26775 701 26776
rect 835 26816 893 26817
rect 835 26776 844 26816
rect 884 26776 893 26816
rect 835 26775 893 26776
rect 19947 26816 19989 26825
rect 19947 26776 19948 26816
rect 19988 26776 19989 26816
rect 19947 26767 19989 26776
rect 20427 26816 20469 26825
rect 20427 26776 20428 26816
rect 20468 26776 20469 26816
rect 20427 26767 20469 26776
rect 20523 26816 20565 26825
rect 20523 26776 20524 26816
rect 20564 26776 20565 26816
rect 20523 26767 20565 26776
rect 20619 26816 20661 26825
rect 20619 26776 20620 26816
rect 20660 26776 20661 26816
rect 20619 26767 20661 26776
rect 29643 26816 29685 26825
rect 29643 26776 29644 26816
rect 29684 26776 29685 26816
rect 29643 26767 29685 26776
rect 30123 26816 30165 26825
rect 30123 26776 30124 26816
rect 30164 26776 30165 26816
rect 30123 26767 30165 26776
rect 34923 26816 34965 26825
rect 34923 26776 34924 26816
rect 34964 26776 34965 26816
rect 34923 26767 34965 26776
rect 35299 26816 35357 26817
rect 35299 26776 35308 26816
rect 35348 26776 35357 26816
rect 35299 26775 35357 26776
rect 36163 26816 36221 26817
rect 36163 26776 36172 26816
rect 36212 26776 36221 26816
rect 36163 26775 36221 26776
rect 20139 26648 20181 26657
rect 20139 26608 20140 26648
rect 20180 26608 20181 26648
rect 20139 26599 20181 26608
rect 20323 26648 20381 26649
rect 20323 26608 20332 26648
rect 20372 26608 20381 26648
rect 20323 26607 20381 26608
rect 576 26480 99360 26504
rect 576 26440 4352 26480
rect 4392 26440 4434 26480
rect 4474 26440 4516 26480
rect 4556 26440 4598 26480
rect 4638 26440 4680 26480
rect 4720 26440 19472 26480
rect 19512 26440 19554 26480
rect 19594 26440 19636 26480
rect 19676 26440 19718 26480
rect 19758 26440 19800 26480
rect 19840 26440 34592 26480
rect 34632 26440 34674 26480
rect 34714 26440 34756 26480
rect 34796 26440 34838 26480
rect 34878 26440 34920 26480
rect 34960 26440 49712 26480
rect 49752 26440 49794 26480
rect 49834 26440 49876 26480
rect 49916 26440 49958 26480
rect 49998 26440 50040 26480
rect 50080 26440 64832 26480
rect 64872 26440 64914 26480
rect 64954 26440 64996 26480
rect 65036 26440 65078 26480
rect 65118 26440 65160 26480
rect 65200 26440 79952 26480
rect 79992 26440 80034 26480
rect 80074 26440 80116 26480
rect 80156 26440 80198 26480
rect 80238 26440 80280 26480
rect 80320 26440 95072 26480
rect 95112 26440 95154 26480
rect 95194 26440 95236 26480
rect 95276 26440 95318 26480
rect 95358 26440 95400 26480
rect 95440 26440 99360 26480
rect 576 26416 99360 26440
rect 17251 26312 17309 26313
rect 17251 26272 17260 26312
rect 17300 26272 17309 26312
rect 17251 26271 17309 26272
rect 21579 26312 21621 26321
rect 21579 26272 21580 26312
rect 21620 26272 21621 26312
rect 21579 26263 21621 26272
rect 25803 26312 25845 26321
rect 25803 26272 25804 26312
rect 25844 26272 25845 26312
rect 25803 26263 25845 26272
rect 28299 26312 28341 26321
rect 28299 26272 28300 26312
rect 28340 26272 28341 26312
rect 28299 26263 28341 26272
rect 14859 26228 14901 26237
rect 14859 26188 14860 26228
rect 14900 26188 14901 26228
rect 14859 26179 14901 26188
rect 643 26144 701 26145
rect 643 26104 652 26144
rect 692 26104 701 26144
rect 643 26103 701 26104
rect 835 26144 893 26145
rect 835 26104 844 26144
rect 884 26104 893 26144
rect 835 26103 893 26104
rect 15235 26144 15293 26145
rect 15235 26104 15244 26144
rect 15284 26104 15293 26144
rect 15235 26103 15293 26104
rect 16099 26144 16157 26145
rect 16099 26104 16108 26144
rect 16148 26104 16157 26144
rect 16099 26103 16157 26104
rect 21483 26144 21525 26153
rect 21483 26104 21484 26144
rect 21524 26104 21525 26144
rect 21483 26095 21525 26104
rect 21675 26144 21717 26153
rect 21675 26104 21676 26144
rect 21716 26104 21717 26144
rect 21675 26095 21717 26104
rect 21771 26144 21813 26153
rect 21771 26104 21772 26144
rect 21812 26104 21813 26144
rect 21771 26095 21813 26104
rect 26379 26144 26421 26153
rect 26379 26104 26380 26144
rect 26420 26104 26421 26144
rect 26379 26095 26421 26104
rect 27235 26144 27293 26145
rect 27235 26104 27244 26144
rect 27284 26104 27293 26144
rect 27235 26103 27293 26104
rect 28299 26144 28341 26153
rect 28299 26104 28300 26144
rect 28340 26104 28341 26144
rect 28299 26095 28341 26104
rect 28387 26144 28445 26145
rect 28387 26104 28396 26144
rect 28436 26104 28445 26144
rect 28387 26103 28445 26104
rect 34339 26144 34397 26145
rect 34339 26104 34348 26144
rect 34388 26104 34397 26144
rect 34339 26103 34397 26104
rect 35299 26144 35357 26145
rect 35299 26104 35308 26144
rect 35348 26104 35357 26144
rect 35299 26103 35357 26104
rect 39619 26144 39677 26145
rect 39619 26104 39628 26144
rect 39668 26104 39677 26144
rect 39619 26103 39677 26104
rect 25987 26060 26045 26061
rect 25987 26020 25996 26060
rect 26036 26020 26045 26060
rect 25987 26019 26045 26020
rect 28203 26060 28245 26069
rect 28203 26020 28204 26060
rect 28244 26020 28245 26060
rect 28203 26011 28245 26020
rect 28107 25976 28149 25985
rect 28107 25936 28108 25976
rect 28148 25936 28149 25976
rect 28107 25927 28149 25936
rect 39915 25892 39957 25901
rect 39915 25852 39916 25892
rect 39956 25852 39957 25892
rect 39915 25843 39957 25852
rect 576 25724 99360 25748
rect 576 25684 3112 25724
rect 3152 25684 3194 25724
rect 3234 25684 3276 25724
rect 3316 25684 3358 25724
rect 3398 25684 3440 25724
rect 3480 25684 18232 25724
rect 18272 25684 18314 25724
rect 18354 25684 18396 25724
rect 18436 25684 18478 25724
rect 18518 25684 18560 25724
rect 18600 25684 33352 25724
rect 33392 25684 33434 25724
rect 33474 25684 33516 25724
rect 33556 25684 33598 25724
rect 33638 25684 33680 25724
rect 33720 25684 48472 25724
rect 48512 25684 48554 25724
rect 48594 25684 48636 25724
rect 48676 25684 48718 25724
rect 48758 25684 48800 25724
rect 48840 25684 63592 25724
rect 63632 25684 63674 25724
rect 63714 25684 63756 25724
rect 63796 25684 63838 25724
rect 63878 25684 63920 25724
rect 63960 25684 78712 25724
rect 78752 25684 78794 25724
rect 78834 25684 78876 25724
rect 78916 25684 78958 25724
rect 78998 25684 79040 25724
rect 79080 25684 93832 25724
rect 93872 25684 93914 25724
rect 93954 25684 93996 25724
rect 94036 25684 94078 25724
rect 94118 25684 94160 25724
rect 94200 25684 99360 25724
rect 576 25660 99360 25684
rect 28195 25556 28253 25557
rect 28195 25516 28204 25556
rect 28244 25516 28253 25556
rect 28195 25515 28253 25516
rect 643 25304 701 25305
rect 643 25264 652 25304
rect 692 25264 701 25304
rect 643 25263 701 25264
rect 835 25304 893 25305
rect 835 25264 844 25304
rect 884 25264 893 25304
rect 835 25263 893 25264
rect 28387 25304 28445 25305
rect 28387 25264 28396 25304
rect 28436 25264 28445 25304
rect 28387 25263 28445 25264
rect 28483 25136 28541 25137
rect 28483 25096 28492 25136
rect 28532 25096 28541 25136
rect 28483 25095 28541 25096
rect 576 24968 99360 24992
rect 576 24928 4352 24968
rect 4392 24928 4434 24968
rect 4474 24928 4516 24968
rect 4556 24928 4598 24968
rect 4638 24928 4680 24968
rect 4720 24928 19472 24968
rect 19512 24928 19554 24968
rect 19594 24928 19636 24968
rect 19676 24928 19718 24968
rect 19758 24928 19800 24968
rect 19840 24928 34592 24968
rect 34632 24928 34674 24968
rect 34714 24928 34756 24968
rect 34796 24928 34838 24968
rect 34878 24928 34920 24968
rect 34960 24928 49712 24968
rect 49752 24928 49794 24968
rect 49834 24928 49876 24968
rect 49916 24928 49958 24968
rect 49998 24928 50040 24968
rect 50080 24928 64832 24968
rect 64872 24928 64914 24968
rect 64954 24928 64996 24968
rect 65036 24928 65078 24968
rect 65118 24928 65160 24968
rect 65200 24928 79952 24968
rect 79992 24928 80034 24968
rect 80074 24928 80116 24968
rect 80156 24928 80198 24968
rect 80238 24928 80280 24968
rect 80320 24928 95072 24968
rect 95112 24928 95154 24968
rect 95194 24928 95236 24968
rect 95276 24928 95318 24968
rect 95358 24928 95400 24968
rect 95440 24928 99360 24968
rect 576 24904 99360 24928
rect 29635 24800 29693 24801
rect 29635 24760 29644 24800
rect 29684 24760 29693 24800
rect 29635 24759 29693 24760
rect 29835 24716 29877 24725
rect 29835 24676 29836 24716
rect 29876 24676 29877 24716
rect 29835 24667 29877 24676
rect 643 24632 701 24633
rect 643 24592 652 24632
rect 692 24592 701 24632
rect 643 24591 701 24592
rect 835 24632 893 24633
rect 835 24592 844 24632
rect 884 24592 893 24632
rect 835 24591 893 24592
rect 23011 24632 23069 24633
rect 23011 24592 23020 24632
rect 23060 24592 23069 24632
rect 23011 24591 23069 24592
rect 23971 24632 24029 24633
rect 23971 24592 23980 24632
rect 24020 24592 24029 24632
rect 23971 24591 24029 24592
rect 30019 24632 30077 24633
rect 30019 24592 30028 24632
rect 30068 24592 30077 24632
rect 30019 24591 30077 24592
rect 22627 24548 22685 24549
rect 22627 24508 22636 24548
rect 22676 24508 22685 24548
rect 22627 24507 22685 24508
rect 576 24212 99360 24236
rect 576 24172 3112 24212
rect 3152 24172 3194 24212
rect 3234 24172 3276 24212
rect 3316 24172 3358 24212
rect 3398 24172 3440 24212
rect 3480 24172 18232 24212
rect 18272 24172 18314 24212
rect 18354 24172 18396 24212
rect 18436 24172 18478 24212
rect 18518 24172 18560 24212
rect 18600 24172 33352 24212
rect 33392 24172 33434 24212
rect 33474 24172 33516 24212
rect 33556 24172 33598 24212
rect 33638 24172 33680 24212
rect 33720 24172 48472 24212
rect 48512 24172 48554 24212
rect 48594 24172 48636 24212
rect 48676 24172 48718 24212
rect 48758 24172 48800 24212
rect 48840 24172 63592 24212
rect 63632 24172 63674 24212
rect 63714 24172 63756 24212
rect 63796 24172 63838 24212
rect 63878 24172 63920 24212
rect 63960 24172 78712 24212
rect 78752 24172 78794 24212
rect 78834 24172 78876 24212
rect 78916 24172 78958 24212
rect 78998 24172 79040 24212
rect 79080 24172 93832 24212
rect 93872 24172 93914 24212
rect 93954 24172 93996 24212
rect 94036 24172 94078 24212
rect 94118 24172 94160 24212
rect 94200 24172 99360 24212
rect 576 24148 99360 24172
rect 28875 23960 28917 23969
rect 28875 23920 28876 23960
rect 28916 23920 28917 23960
rect 28875 23911 28917 23920
rect 32803 23876 32861 23877
rect 32803 23836 32812 23876
rect 32852 23836 32861 23876
rect 32803 23835 32861 23836
rect 643 23792 701 23793
rect 643 23752 652 23792
rect 692 23752 701 23792
rect 643 23751 701 23752
rect 835 23792 893 23793
rect 835 23752 844 23792
rect 884 23752 893 23792
rect 835 23751 893 23752
rect 28963 23792 29021 23793
rect 28963 23752 28972 23792
rect 29012 23752 29021 23792
rect 28963 23751 29021 23752
rect 33283 23792 33341 23793
rect 33283 23752 33292 23792
rect 33332 23752 33341 23792
rect 33283 23751 33341 23752
rect 33771 23624 33813 23633
rect 33771 23584 33772 23624
rect 33812 23584 33813 23624
rect 33771 23575 33813 23584
rect 576 23456 99360 23480
rect 576 23416 4352 23456
rect 4392 23416 4434 23456
rect 4474 23416 4516 23456
rect 4556 23416 4598 23456
rect 4638 23416 4680 23456
rect 4720 23416 19472 23456
rect 19512 23416 19554 23456
rect 19594 23416 19636 23456
rect 19676 23416 19718 23456
rect 19758 23416 19800 23456
rect 19840 23416 34592 23456
rect 34632 23416 34674 23456
rect 34714 23416 34756 23456
rect 34796 23416 34838 23456
rect 34878 23416 34920 23456
rect 34960 23416 49712 23456
rect 49752 23416 49794 23456
rect 49834 23416 49876 23456
rect 49916 23416 49958 23456
rect 49998 23416 50040 23456
rect 50080 23416 64832 23456
rect 64872 23416 64914 23456
rect 64954 23416 64996 23456
rect 65036 23416 65078 23456
rect 65118 23416 65160 23456
rect 65200 23416 79952 23456
rect 79992 23416 80034 23456
rect 80074 23416 80116 23456
rect 80156 23416 80198 23456
rect 80238 23416 80280 23456
rect 80320 23416 95072 23456
rect 95112 23416 95154 23456
rect 95194 23416 95236 23456
rect 95276 23416 95318 23456
rect 95358 23416 95400 23456
rect 95440 23416 99360 23456
rect 576 23392 99360 23416
rect 19371 23120 19413 23129
rect 19371 23080 19372 23120
rect 19412 23080 19413 23120
rect 19371 23071 19413 23080
rect 19747 23120 19805 23121
rect 19747 23080 19756 23120
rect 19796 23080 19805 23120
rect 19747 23079 19805 23080
rect 20611 23120 20669 23121
rect 20611 23080 20620 23120
rect 20660 23080 20669 23120
rect 20611 23079 20669 23080
rect 28579 23120 28637 23121
rect 28579 23080 28588 23120
rect 28628 23080 28637 23120
rect 28579 23079 28637 23080
rect 28683 23120 28725 23129
rect 28683 23080 28684 23120
rect 28724 23080 28725 23120
rect 28683 23071 28725 23080
rect 28867 23120 28925 23121
rect 28867 23080 28876 23120
rect 28916 23080 28925 23120
rect 28867 23079 28925 23080
rect 34059 23120 34101 23129
rect 34059 23080 34060 23120
rect 34100 23080 34101 23120
rect 34059 23071 34101 23080
rect 34435 23120 34493 23121
rect 34435 23080 34444 23120
rect 34484 23080 34493 23120
rect 34435 23079 34493 23080
rect 35299 23120 35357 23121
rect 35299 23080 35308 23120
rect 35348 23080 35357 23120
rect 35299 23079 35357 23080
rect 21763 22868 21821 22869
rect 21763 22828 21772 22868
rect 21812 22828 21821 22868
rect 21763 22827 21821 22828
rect 28875 22868 28917 22877
rect 28875 22828 28876 22868
rect 28916 22828 28917 22868
rect 28875 22819 28917 22828
rect 36451 22868 36509 22869
rect 36451 22828 36460 22868
rect 36500 22828 36509 22868
rect 36451 22827 36509 22828
rect 576 22700 99360 22724
rect 576 22660 3112 22700
rect 3152 22660 3194 22700
rect 3234 22660 3276 22700
rect 3316 22660 3358 22700
rect 3398 22660 3440 22700
rect 3480 22660 18232 22700
rect 18272 22660 18314 22700
rect 18354 22660 18396 22700
rect 18436 22660 18478 22700
rect 18518 22660 18560 22700
rect 18600 22660 33352 22700
rect 33392 22660 33434 22700
rect 33474 22660 33516 22700
rect 33556 22660 33598 22700
rect 33638 22660 33680 22700
rect 33720 22660 48472 22700
rect 48512 22660 48554 22700
rect 48594 22660 48636 22700
rect 48676 22660 48718 22700
rect 48758 22660 48800 22700
rect 48840 22660 63592 22700
rect 63632 22660 63674 22700
rect 63714 22660 63756 22700
rect 63796 22660 63838 22700
rect 63878 22660 63920 22700
rect 63960 22660 78712 22700
rect 78752 22660 78794 22700
rect 78834 22660 78876 22700
rect 78916 22660 78958 22700
rect 78998 22660 79040 22700
rect 79080 22660 93832 22700
rect 93872 22660 93914 22700
rect 93954 22660 93996 22700
rect 94036 22660 94078 22700
rect 94118 22660 94160 22700
rect 94200 22660 99360 22700
rect 576 22636 99360 22660
rect 651 22448 693 22457
rect 651 22408 652 22448
rect 692 22408 693 22448
rect 651 22399 693 22408
rect 29163 22448 29205 22457
rect 29163 22408 29164 22448
rect 29204 22408 29205 22448
rect 29163 22399 29205 22408
rect 26571 22364 26613 22373
rect 26571 22324 26572 22364
rect 26612 22324 26613 22364
rect 26571 22315 26613 22324
rect 35307 22364 35349 22373
rect 35307 22324 35308 22364
rect 35348 22324 35349 22364
rect 35307 22315 35349 22324
rect 41547 22364 41589 22373
rect 41547 22324 41548 22364
rect 41588 22324 41589 22364
rect 41547 22315 41589 22324
rect 15331 22280 15389 22281
rect 15331 22240 15340 22280
rect 15380 22240 15389 22280
rect 15331 22239 15389 22240
rect 16195 22280 16253 22281
rect 16195 22240 16204 22280
rect 16244 22240 16253 22280
rect 16195 22239 16253 22240
rect 24547 22280 24605 22281
rect 24547 22240 24556 22280
rect 24596 22240 24605 22280
rect 24547 22239 24605 22240
rect 25411 22280 25469 22281
rect 25411 22240 25420 22280
rect 25460 22240 25469 22280
rect 25411 22239 25469 22240
rect 28683 22280 28725 22289
rect 28683 22240 28684 22280
rect 28724 22240 28725 22280
rect 28683 22231 28725 22240
rect 28779 22280 28821 22289
rect 28779 22240 28780 22280
rect 28820 22240 28821 22280
rect 28779 22231 28821 22240
rect 28875 22280 28917 22289
rect 28875 22240 28876 22280
rect 28916 22240 28917 22280
rect 28875 22231 28917 22240
rect 29251 22280 29309 22281
rect 29251 22240 29260 22280
rect 29300 22240 29309 22280
rect 29251 22239 29309 22240
rect 32419 22280 32477 22281
rect 32419 22240 32428 22280
rect 32468 22240 32477 22280
rect 32419 22239 32477 22240
rect 32523 22280 32565 22289
rect 32523 22240 32524 22280
rect 32564 22240 32565 22280
rect 32523 22231 32565 22240
rect 32619 22280 32661 22289
rect 32619 22240 32620 22280
rect 32660 22240 32661 22280
rect 32619 22231 32661 22240
rect 34059 22280 34101 22289
rect 34059 22240 34060 22280
rect 34100 22240 34101 22280
rect 34059 22231 34101 22240
rect 34155 22280 34197 22289
rect 34155 22240 34156 22280
rect 34196 22240 34197 22280
rect 34155 22231 34197 22240
rect 34923 22280 34965 22289
rect 34923 22240 34924 22280
rect 34964 22240 34965 22280
rect 34923 22231 34965 22240
rect 35019 22280 35061 22289
rect 35019 22240 35020 22280
rect 35060 22240 35061 22280
rect 35019 22231 35061 22240
rect 35211 22280 35253 22289
rect 35211 22240 35212 22280
rect 35252 22240 35253 22280
rect 35211 22231 35253 22240
rect 35395 22280 35453 22281
rect 35395 22240 35404 22280
rect 35444 22240 35453 22280
rect 35395 22239 35453 22240
rect 35595 22280 35637 22289
rect 35595 22240 35596 22280
rect 35636 22240 35637 22280
rect 35595 22231 35637 22240
rect 35779 22280 35837 22281
rect 35779 22240 35788 22280
rect 35828 22240 35837 22280
rect 35779 22239 35837 22240
rect 39523 22280 39581 22281
rect 39523 22240 39532 22280
rect 39572 22240 39581 22280
rect 39523 22239 39581 22240
rect 40387 22280 40445 22281
rect 40387 22240 40396 22280
rect 40436 22240 40445 22280
rect 40387 22239 40445 22240
rect 14955 22196 14997 22205
rect 14955 22156 14956 22196
rect 14996 22156 14997 22196
rect 14955 22147 14997 22156
rect 24171 22196 24213 22205
rect 24171 22156 24172 22196
rect 24212 22156 24213 22196
rect 24171 22147 24213 22156
rect 34243 22196 34301 22197
rect 34243 22156 34252 22196
rect 34292 22156 34301 22196
rect 34243 22155 34301 22156
rect 34811 22196 34869 22197
rect 34811 22156 34820 22196
rect 34860 22156 34869 22196
rect 34811 22155 34869 22156
rect 35691 22196 35733 22205
rect 35691 22156 35692 22196
rect 35732 22156 35733 22196
rect 35691 22147 35733 22156
rect 39147 22196 39189 22205
rect 39147 22156 39148 22196
rect 39188 22156 39189 22196
rect 39147 22147 39189 22156
rect 17347 22112 17405 22113
rect 17347 22072 17356 22112
rect 17396 22072 17405 22112
rect 17347 22071 17405 22072
rect 28963 22112 29021 22113
rect 28963 22072 28972 22112
rect 29012 22072 29021 22112
rect 28963 22071 29021 22072
rect 34339 22112 34397 22113
rect 34339 22072 34348 22112
rect 34388 22072 34397 22112
rect 34339 22071 34397 22072
rect 34443 22112 34485 22121
rect 34443 22072 34444 22112
rect 34484 22072 34485 22112
rect 34443 22063 34485 22072
rect 34635 22112 34677 22121
rect 34635 22072 34636 22112
rect 34676 22072 34677 22112
rect 34635 22063 34677 22072
rect 34723 22112 34781 22113
rect 34723 22072 34732 22112
rect 34772 22072 34781 22112
rect 34723 22071 34781 22072
rect 576 21944 99360 21968
rect 576 21904 4352 21944
rect 4392 21904 4434 21944
rect 4474 21904 4516 21944
rect 4556 21904 4598 21944
rect 4638 21904 4680 21944
rect 4720 21904 19472 21944
rect 19512 21904 19554 21944
rect 19594 21904 19636 21944
rect 19676 21904 19718 21944
rect 19758 21904 19800 21944
rect 19840 21904 34592 21944
rect 34632 21904 34674 21944
rect 34714 21904 34756 21944
rect 34796 21904 34838 21944
rect 34878 21904 34920 21944
rect 34960 21904 49712 21944
rect 49752 21904 49794 21944
rect 49834 21904 49876 21944
rect 49916 21904 49958 21944
rect 49998 21904 50040 21944
rect 50080 21904 64832 21944
rect 64872 21904 64914 21944
rect 64954 21904 64996 21944
rect 65036 21904 65078 21944
rect 65118 21904 65160 21944
rect 65200 21904 79952 21944
rect 79992 21904 80034 21944
rect 80074 21904 80116 21944
rect 80156 21904 80198 21944
rect 80238 21904 80280 21944
rect 80320 21904 95072 21944
rect 95112 21904 95154 21944
rect 95194 21904 95236 21944
rect 95276 21904 95318 21944
rect 95358 21904 95400 21944
rect 95440 21904 99360 21944
rect 576 21880 99360 21904
rect 28387 21608 28445 21609
rect 28387 21568 28396 21608
rect 28436 21568 28445 21608
rect 28387 21567 28445 21568
rect 29347 21608 29405 21609
rect 29347 21568 29356 21608
rect 29396 21568 29405 21608
rect 29347 21567 29405 21568
rect 576 21188 99360 21212
rect 576 21148 3112 21188
rect 3152 21148 3194 21188
rect 3234 21148 3276 21188
rect 3316 21148 3358 21188
rect 3398 21148 3440 21188
rect 3480 21148 18232 21188
rect 18272 21148 18314 21188
rect 18354 21148 18396 21188
rect 18436 21148 18478 21188
rect 18518 21148 18560 21188
rect 18600 21148 33352 21188
rect 33392 21148 33434 21188
rect 33474 21148 33516 21188
rect 33556 21148 33598 21188
rect 33638 21148 33680 21188
rect 33720 21148 48472 21188
rect 48512 21148 48554 21188
rect 48594 21148 48636 21188
rect 48676 21148 48718 21188
rect 48758 21148 48800 21188
rect 48840 21148 63592 21188
rect 63632 21148 63674 21188
rect 63714 21148 63756 21188
rect 63796 21148 63838 21188
rect 63878 21148 63920 21188
rect 63960 21148 78712 21188
rect 78752 21148 78794 21188
rect 78834 21148 78876 21188
rect 78916 21148 78958 21188
rect 78998 21148 79040 21188
rect 79080 21148 93832 21188
rect 93872 21148 93914 21188
rect 93954 21148 93996 21188
rect 94036 21148 94078 21188
rect 94118 21148 94160 21188
rect 94200 21148 99360 21188
rect 576 21124 99360 21148
rect 19171 21020 19229 21021
rect 19171 20980 19180 21020
rect 19220 20980 19229 21020
rect 19171 20979 19229 20980
rect 651 20936 693 20945
rect 651 20896 652 20936
rect 692 20896 693 20936
rect 651 20887 693 20896
rect 30595 20936 30653 20937
rect 30595 20896 30604 20936
rect 30644 20896 30653 20936
rect 30595 20895 30653 20896
rect 30795 20852 30837 20861
rect 30795 20812 30796 20852
rect 30836 20812 30837 20852
rect 30795 20803 30837 20812
rect 31363 20852 31421 20853
rect 31363 20812 31372 20852
rect 31412 20812 31421 20852
rect 31363 20811 31421 20812
rect 19371 20768 19413 20777
rect 19371 20728 19372 20768
rect 19412 20728 19413 20768
rect 19371 20719 19413 20728
rect 19467 20768 19509 20777
rect 19467 20728 19468 20768
rect 19508 20728 19509 20768
rect 19467 20719 19509 20728
rect 19563 20768 19605 20777
rect 19563 20728 19564 20768
rect 19604 20728 19605 20768
rect 19563 20719 19605 20728
rect 22635 20768 22677 20777
rect 22635 20728 22636 20768
rect 22676 20728 22677 20768
rect 22635 20719 22677 20728
rect 22731 20768 22773 20777
rect 22731 20728 22732 20768
rect 22772 20728 22773 20768
rect 22731 20719 22773 20728
rect 22827 20768 22869 20777
rect 22827 20728 22828 20768
rect 22868 20728 22869 20768
rect 22827 20719 22869 20728
rect 23115 20768 23157 20777
rect 23115 20728 23116 20768
rect 23156 20728 23157 20768
rect 23115 20719 23157 20728
rect 23211 20768 23253 20777
rect 23211 20728 23212 20768
rect 23252 20728 23253 20768
rect 23211 20719 23253 20728
rect 23307 20768 23349 20777
rect 23307 20728 23308 20768
rect 23348 20728 23349 20768
rect 23307 20719 23349 20728
rect 23403 20768 23445 20777
rect 23403 20728 23404 20768
rect 23444 20728 23445 20768
rect 23403 20719 23445 20728
rect 29163 20768 29205 20777
rect 29163 20728 29164 20768
rect 29204 20728 29205 20768
rect 29163 20719 29205 20728
rect 30315 20768 30357 20777
rect 30315 20728 30316 20768
rect 30356 20728 30357 20768
rect 30315 20719 30357 20728
rect 30507 20768 30549 20777
rect 30507 20728 30508 20768
rect 30548 20728 30549 20768
rect 30507 20719 30549 20728
rect 30603 20768 30645 20777
rect 30603 20728 30604 20768
rect 30644 20728 30645 20768
rect 30603 20719 30645 20728
rect 31171 20768 31229 20769
rect 31171 20728 31180 20768
rect 31220 20728 31229 20768
rect 31171 20727 31229 20728
rect 22923 20684 22965 20693
rect 22923 20644 22924 20684
rect 22964 20644 22965 20684
rect 22923 20635 22965 20644
rect 29443 20600 29501 20601
rect 29443 20560 29452 20600
rect 29492 20560 29501 20600
rect 29443 20559 29501 20560
rect 29635 20600 29693 20601
rect 29635 20560 29644 20600
rect 29684 20560 29693 20600
rect 29635 20559 29693 20560
rect 30883 20600 30941 20601
rect 30883 20560 30892 20600
rect 30932 20560 30941 20600
rect 30883 20559 30941 20560
rect 576 20432 99360 20456
rect 576 20392 4352 20432
rect 4392 20392 4434 20432
rect 4474 20392 4516 20432
rect 4556 20392 4598 20432
rect 4638 20392 4680 20432
rect 4720 20392 19472 20432
rect 19512 20392 19554 20432
rect 19594 20392 19636 20432
rect 19676 20392 19718 20432
rect 19758 20392 19800 20432
rect 19840 20392 34592 20432
rect 34632 20392 34674 20432
rect 34714 20392 34756 20432
rect 34796 20392 34838 20432
rect 34878 20392 34920 20432
rect 34960 20392 49712 20432
rect 49752 20392 49794 20432
rect 49834 20392 49876 20432
rect 49916 20392 49958 20432
rect 49998 20392 50040 20432
rect 50080 20392 64832 20432
rect 64872 20392 64914 20432
rect 64954 20392 64996 20432
rect 65036 20392 65078 20432
rect 65118 20392 65160 20432
rect 65200 20392 79952 20432
rect 79992 20392 80034 20432
rect 80074 20392 80116 20432
rect 80156 20392 80198 20432
rect 80238 20392 80280 20432
rect 80320 20392 95072 20432
rect 95112 20392 95154 20432
rect 95194 20392 95236 20432
rect 95276 20392 95318 20432
rect 95358 20392 95400 20432
rect 95440 20392 99360 20432
rect 576 20368 99360 20392
rect 22051 20264 22109 20265
rect 22051 20224 22060 20264
rect 22100 20224 22109 20264
rect 22051 20223 22109 20224
rect 15427 20180 15485 20181
rect 15427 20140 15436 20180
rect 15476 20140 15485 20180
rect 15427 20139 15485 20140
rect 34923 20180 34965 20189
rect 34923 20140 34924 20180
rect 34964 20140 34965 20180
rect 34923 20131 34965 20140
rect 15619 20096 15677 20097
rect 15619 20056 15628 20096
rect 15668 20056 15677 20096
rect 15619 20055 15677 20056
rect 15907 20096 15965 20097
rect 15907 20056 15916 20096
rect 15956 20056 15965 20096
rect 15907 20055 15965 20056
rect 21091 20096 21149 20097
rect 21091 20056 21100 20096
rect 21140 20056 21149 20096
rect 21091 20055 21149 20056
rect 21195 20096 21237 20105
rect 21195 20056 21196 20096
rect 21236 20056 21237 20096
rect 21195 20047 21237 20056
rect 21379 20096 21437 20097
rect 21379 20056 21388 20096
rect 21428 20056 21437 20096
rect 21379 20055 21437 20056
rect 21771 20096 21813 20105
rect 21771 20056 21772 20096
rect 21812 20056 21813 20096
rect 21771 20047 21813 20056
rect 21867 20096 21909 20105
rect 21867 20056 21868 20096
rect 21908 20056 21909 20096
rect 21867 20047 21909 20056
rect 23203 20096 23261 20097
rect 23203 20056 23212 20096
rect 23252 20056 23261 20096
rect 23203 20055 23261 20056
rect 24163 20096 24221 20097
rect 24163 20056 24172 20096
rect 24212 20056 24221 20096
rect 24163 20055 24221 20056
rect 34827 20096 34869 20105
rect 34827 20056 34828 20096
rect 34868 20056 34869 20096
rect 34827 20047 34869 20056
rect 35011 20096 35069 20097
rect 35011 20056 35020 20096
rect 35060 20056 35069 20096
rect 35011 20055 35069 20056
rect 39907 20096 39965 20097
rect 39907 20056 39916 20096
rect 39956 20056 39965 20096
rect 39907 20055 39965 20056
rect 22819 20012 22877 20013
rect 22819 19972 22828 20012
rect 22868 19972 22877 20012
rect 22819 19971 22877 19972
rect 651 19928 693 19937
rect 651 19888 652 19928
rect 692 19888 693 19928
rect 651 19879 693 19888
rect 21387 19928 21429 19937
rect 21387 19888 21388 19928
rect 21428 19888 21429 19928
rect 21387 19879 21429 19888
rect 23691 19844 23733 19853
rect 23691 19804 23692 19844
rect 23732 19804 23733 19844
rect 23691 19795 23733 19804
rect 39235 19844 39293 19845
rect 39235 19804 39244 19844
rect 39284 19804 39293 19844
rect 39235 19803 39293 19804
rect 576 19676 99360 19700
rect 576 19636 3112 19676
rect 3152 19636 3194 19676
rect 3234 19636 3276 19676
rect 3316 19636 3358 19676
rect 3398 19636 3440 19676
rect 3480 19636 18232 19676
rect 18272 19636 18314 19676
rect 18354 19636 18396 19676
rect 18436 19636 18478 19676
rect 18518 19636 18560 19676
rect 18600 19636 33352 19676
rect 33392 19636 33434 19676
rect 33474 19636 33516 19676
rect 33556 19636 33598 19676
rect 33638 19636 33680 19676
rect 33720 19636 48472 19676
rect 48512 19636 48554 19676
rect 48594 19636 48636 19676
rect 48676 19636 48718 19676
rect 48758 19636 48800 19676
rect 48840 19636 63592 19676
rect 63632 19636 63674 19676
rect 63714 19636 63756 19676
rect 63796 19636 63838 19676
rect 63878 19636 63920 19676
rect 63960 19636 78712 19676
rect 78752 19636 78794 19676
rect 78834 19636 78876 19676
rect 78916 19636 78958 19676
rect 78998 19636 79040 19676
rect 79080 19636 93832 19676
rect 93872 19636 93914 19676
rect 93954 19636 93996 19676
rect 94036 19636 94078 19676
rect 94118 19636 94160 19676
rect 94200 19636 99360 19676
rect 576 19612 99360 19636
rect 41155 19508 41213 19509
rect 41155 19468 41164 19508
rect 41204 19468 41213 19508
rect 41155 19467 41213 19468
rect 651 19424 693 19433
rect 651 19384 652 19424
rect 692 19384 693 19424
rect 651 19375 693 19384
rect 33867 19424 33909 19433
rect 33867 19384 33868 19424
rect 33908 19384 33909 19424
rect 33867 19375 33909 19384
rect 37507 19424 37565 19425
rect 37507 19384 37516 19424
rect 37556 19384 37565 19424
rect 37507 19383 37565 19384
rect 19179 19340 19221 19349
rect 19179 19300 19180 19340
rect 19220 19300 19221 19340
rect 19179 19291 19221 19300
rect 19083 19256 19125 19265
rect 19083 19216 19084 19256
rect 19124 19216 19125 19256
rect 19083 19207 19125 19216
rect 19459 19256 19517 19257
rect 19459 19216 19468 19256
rect 19508 19216 19517 19256
rect 19459 19215 19517 19216
rect 19651 19256 19709 19257
rect 19651 19216 19660 19256
rect 19700 19216 19709 19256
rect 19651 19215 19709 19216
rect 33187 19256 33245 19257
rect 33187 19216 33196 19256
rect 33236 19216 33245 19256
rect 33187 19215 33245 19216
rect 36835 19256 36893 19257
rect 36835 19216 36844 19256
rect 36884 19216 36893 19256
rect 36835 19215 36893 19216
rect 37131 19256 37173 19265
rect 37131 19216 37132 19256
rect 37172 19216 37173 19256
rect 37131 19207 37173 19216
rect 37227 19256 37269 19265
rect 37227 19216 37228 19256
rect 37268 19216 37269 19256
rect 37227 19207 37269 19216
rect 38763 19256 38805 19265
rect 38763 19216 38764 19256
rect 38804 19216 38805 19256
rect 38763 19207 38805 19216
rect 39139 19256 39197 19257
rect 39139 19216 39148 19256
rect 39188 19216 39197 19256
rect 39139 19215 39197 19216
rect 40003 19256 40061 19257
rect 40003 19216 40012 19256
rect 40052 19216 40061 19256
rect 40003 19215 40061 19216
rect 19467 19088 19509 19097
rect 19467 19048 19468 19088
rect 19508 19048 19509 19088
rect 19467 19039 19509 19048
rect 576 18920 99360 18944
rect 576 18880 4352 18920
rect 4392 18880 4434 18920
rect 4474 18880 4516 18920
rect 4556 18880 4598 18920
rect 4638 18880 4680 18920
rect 4720 18880 19472 18920
rect 19512 18880 19554 18920
rect 19594 18880 19636 18920
rect 19676 18880 19718 18920
rect 19758 18880 19800 18920
rect 19840 18880 34592 18920
rect 34632 18880 34674 18920
rect 34714 18880 34756 18920
rect 34796 18880 34838 18920
rect 34878 18880 34920 18920
rect 34960 18880 49712 18920
rect 49752 18880 49794 18920
rect 49834 18880 49876 18920
rect 49916 18880 49958 18920
rect 49998 18880 50040 18920
rect 50080 18880 64832 18920
rect 64872 18880 64914 18920
rect 64954 18880 64996 18920
rect 65036 18880 65078 18920
rect 65118 18880 65160 18920
rect 65200 18880 79952 18920
rect 79992 18880 80034 18920
rect 80074 18880 80116 18920
rect 80156 18880 80198 18920
rect 80238 18880 80280 18920
rect 80320 18880 95072 18920
rect 95112 18880 95154 18920
rect 95194 18880 95236 18920
rect 95276 18880 95318 18920
rect 95358 18880 95400 18920
rect 95440 18880 99360 18920
rect 576 18856 99360 18880
rect 17539 18668 17597 18669
rect 17539 18628 17548 18668
rect 17588 18628 17597 18668
rect 17539 18627 17597 18628
rect 27339 18668 27381 18677
rect 27339 18628 27340 18668
rect 27380 18628 27381 18668
rect 27339 18619 27381 18628
rect 17731 18584 17789 18585
rect 17731 18544 17740 18584
rect 17780 18544 17789 18584
rect 17731 18543 17789 18544
rect 18019 18584 18077 18585
rect 18019 18544 18028 18584
rect 18068 18544 18077 18584
rect 18019 18543 18077 18544
rect 22443 18584 22485 18593
rect 22443 18544 22444 18584
rect 22484 18544 22485 18584
rect 22443 18535 22485 18544
rect 26083 18584 26141 18585
rect 26083 18544 26092 18584
rect 26132 18544 26141 18584
rect 26083 18543 26141 18544
rect 26475 18584 26517 18593
rect 26475 18544 26476 18584
rect 26516 18544 26517 18584
rect 26475 18535 26517 18544
rect 27427 18584 27485 18585
rect 27427 18544 27436 18584
rect 27476 18544 27485 18584
rect 27427 18543 27485 18544
rect 28395 18584 28437 18593
rect 28395 18544 28396 18584
rect 28436 18544 28437 18584
rect 28395 18535 28437 18544
rect 29059 18584 29117 18585
rect 29059 18544 29068 18584
rect 29108 18544 29117 18584
rect 29059 18543 29117 18544
rect 22251 18500 22293 18509
rect 22251 18460 22252 18500
rect 22292 18460 22293 18500
rect 22251 18451 22293 18460
rect 26187 18500 26229 18509
rect 26187 18460 26188 18500
rect 26228 18460 26229 18500
rect 26187 18451 26229 18460
rect 26379 18500 26421 18509
rect 26379 18460 26380 18500
rect 26420 18460 26421 18500
rect 26379 18451 26421 18460
rect 651 18416 693 18425
rect 651 18376 652 18416
rect 692 18376 693 18416
rect 651 18367 693 18376
rect 26283 18416 26325 18425
rect 26283 18376 26284 18416
rect 26324 18376 26325 18416
rect 26283 18367 26325 18376
rect 22443 18332 22485 18341
rect 22443 18292 22444 18332
rect 22484 18292 22485 18332
rect 22443 18283 22485 18292
rect 576 18164 99360 18188
rect 576 18124 3112 18164
rect 3152 18124 3194 18164
rect 3234 18124 3276 18164
rect 3316 18124 3358 18164
rect 3398 18124 3440 18164
rect 3480 18124 18232 18164
rect 18272 18124 18314 18164
rect 18354 18124 18396 18164
rect 18436 18124 18478 18164
rect 18518 18124 18560 18164
rect 18600 18124 33352 18164
rect 33392 18124 33434 18164
rect 33474 18124 33516 18164
rect 33556 18124 33598 18164
rect 33638 18124 33680 18164
rect 33720 18124 48472 18164
rect 48512 18124 48554 18164
rect 48594 18124 48636 18164
rect 48676 18124 48718 18164
rect 48758 18124 48800 18164
rect 48840 18124 63592 18164
rect 63632 18124 63674 18164
rect 63714 18124 63756 18164
rect 63796 18124 63838 18164
rect 63878 18124 63920 18164
rect 63960 18124 78712 18164
rect 78752 18124 78794 18164
rect 78834 18124 78876 18164
rect 78916 18124 78958 18164
rect 78998 18124 79040 18164
rect 79080 18124 93832 18164
rect 93872 18124 93914 18164
rect 93954 18124 93996 18164
rect 94036 18124 94078 18164
rect 94118 18124 94160 18164
rect 94200 18124 99360 18164
rect 576 18100 99360 18124
rect 21387 17996 21429 18005
rect 21387 17956 21388 17996
rect 21428 17956 21429 17996
rect 21387 17947 21429 17956
rect 21867 17996 21909 18005
rect 21867 17956 21868 17996
rect 21908 17956 21909 17996
rect 21867 17947 21909 17956
rect 651 17912 693 17921
rect 651 17872 652 17912
rect 692 17872 693 17912
rect 651 17863 693 17872
rect 22819 17912 22877 17913
rect 22819 17872 22828 17912
rect 22868 17872 22877 17912
rect 22819 17871 22877 17872
rect 29163 17828 29205 17837
rect 29163 17788 29164 17828
rect 29204 17788 29205 17828
rect 29163 17779 29205 17788
rect 16099 17744 16157 17745
rect 16099 17704 16108 17744
rect 16148 17704 16157 17744
rect 16099 17703 16157 17704
rect 16203 17744 16245 17753
rect 16203 17704 16204 17744
rect 16244 17704 16245 17744
rect 16203 17695 16245 17704
rect 21283 17744 21341 17745
rect 21283 17704 21292 17744
rect 21332 17704 21341 17744
rect 21283 17703 21341 17704
rect 21763 17744 21821 17745
rect 21763 17704 21772 17744
rect 21812 17704 21821 17744
rect 21763 17703 21821 17704
rect 22155 17744 22197 17753
rect 22155 17704 22156 17744
rect 22196 17704 22197 17744
rect 22155 17695 22197 17704
rect 22347 17744 22389 17753
rect 22347 17704 22348 17744
rect 22388 17704 22389 17744
rect 22347 17695 22389 17704
rect 22539 17744 22581 17753
rect 22539 17704 22540 17744
rect 22580 17704 22581 17744
rect 22539 17695 22581 17704
rect 22731 17744 22773 17753
rect 22731 17704 22732 17744
rect 22772 17704 22773 17744
rect 22731 17695 22773 17704
rect 22827 17744 22869 17753
rect 22827 17704 22828 17744
rect 22868 17704 22869 17744
rect 22827 17695 22869 17704
rect 26763 17744 26805 17753
rect 26763 17704 26764 17744
rect 26804 17704 26805 17744
rect 26763 17695 26805 17704
rect 27139 17744 27197 17745
rect 27139 17704 27148 17744
rect 27188 17704 27197 17744
rect 27139 17703 27197 17704
rect 28003 17744 28061 17745
rect 28003 17704 28012 17744
rect 28052 17704 28061 17744
rect 28003 17703 28061 17704
rect 33675 17744 33717 17753
rect 33675 17704 33676 17744
rect 33716 17704 33717 17744
rect 33675 17695 33717 17704
rect 33859 17744 33917 17745
rect 33859 17704 33868 17744
rect 33908 17704 33917 17744
rect 33859 17703 33917 17704
rect 37891 17744 37949 17745
rect 37891 17704 37900 17744
rect 37940 17704 37949 17744
rect 37891 17703 37949 17704
rect 38763 17744 38805 17753
rect 38763 17704 38764 17744
rect 38804 17704 38805 17744
rect 38763 17695 38805 17704
rect 22251 17660 22293 17669
rect 22251 17620 22252 17660
rect 22292 17620 22293 17660
rect 22251 17611 22293 17620
rect 33771 17660 33813 17669
rect 33771 17620 33772 17660
rect 33812 17620 33813 17660
rect 33771 17611 33813 17620
rect 15819 17576 15861 17585
rect 15819 17536 15820 17576
rect 15860 17536 15861 17576
rect 15819 17527 15861 17536
rect 576 17408 99360 17432
rect 576 17368 4352 17408
rect 4392 17368 4434 17408
rect 4474 17368 4516 17408
rect 4556 17368 4598 17408
rect 4638 17368 4680 17408
rect 4720 17368 19472 17408
rect 19512 17368 19554 17408
rect 19594 17368 19636 17408
rect 19676 17368 19718 17408
rect 19758 17368 19800 17408
rect 19840 17368 34592 17408
rect 34632 17368 34674 17408
rect 34714 17368 34756 17408
rect 34796 17368 34838 17408
rect 34878 17368 34920 17408
rect 34960 17368 49712 17408
rect 49752 17368 49794 17408
rect 49834 17368 49876 17408
rect 49916 17368 49958 17408
rect 49998 17368 50040 17408
rect 50080 17368 64832 17408
rect 64872 17368 64914 17408
rect 64954 17368 64996 17408
rect 65036 17368 65078 17408
rect 65118 17368 65160 17408
rect 65200 17368 79952 17408
rect 79992 17368 80034 17408
rect 80074 17368 80116 17408
rect 80156 17368 80198 17408
rect 80238 17368 80280 17408
rect 80320 17368 95072 17408
rect 95112 17368 95154 17408
rect 95194 17368 95236 17408
rect 95276 17368 95318 17408
rect 95358 17368 95400 17408
rect 95440 17368 99360 17408
rect 576 17344 99360 17368
rect 31371 17156 31413 17165
rect 31371 17116 31372 17156
rect 31412 17116 31413 17156
rect 31371 17107 31413 17116
rect 15819 17072 15861 17081
rect 15819 17032 15820 17072
rect 15860 17032 15861 17072
rect 15819 17023 15861 17032
rect 16011 17072 16053 17081
rect 16011 17032 16012 17072
rect 16052 17032 16053 17072
rect 16011 17023 16053 17032
rect 22059 17072 22101 17081
rect 22059 17032 22060 17072
rect 22100 17032 22101 17072
rect 22059 17023 22101 17032
rect 22251 17072 22293 17081
rect 22251 17032 22252 17072
rect 22292 17032 22293 17072
rect 22251 17023 22293 17032
rect 22347 17072 22389 17081
rect 22347 17032 22348 17072
rect 22388 17032 22389 17072
rect 22347 17023 22389 17032
rect 31747 17072 31805 17073
rect 31747 17032 31756 17072
rect 31796 17032 31805 17072
rect 31747 17031 31805 17032
rect 32611 17072 32669 17073
rect 32611 17032 32620 17072
rect 32660 17032 32669 17072
rect 32611 17031 32669 17032
rect 34251 17072 34293 17081
rect 34251 17032 34252 17072
rect 34292 17032 34293 17072
rect 34251 17023 34293 17032
rect 15915 16988 15957 16997
rect 15915 16948 15916 16988
rect 15956 16948 15957 16988
rect 15915 16939 15957 16948
rect 33771 16988 33813 16997
rect 33771 16948 33772 16988
rect 33812 16948 33813 16988
rect 33771 16939 33813 16948
rect 34059 16988 34101 16997
rect 34059 16948 34060 16988
rect 34100 16948 34101 16988
rect 34059 16939 34101 16948
rect 651 16904 693 16913
rect 651 16864 652 16904
rect 692 16864 693 16904
rect 651 16855 693 16864
rect 22339 16904 22397 16905
rect 22339 16864 22348 16904
rect 22388 16864 22397 16904
rect 22339 16863 22397 16864
rect 34251 16820 34293 16829
rect 34251 16780 34252 16820
rect 34292 16780 34293 16820
rect 34251 16771 34293 16780
rect 576 16652 99360 16676
rect 576 16612 3112 16652
rect 3152 16612 3194 16652
rect 3234 16612 3276 16652
rect 3316 16612 3358 16652
rect 3398 16612 3440 16652
rect 3480 16612 18232 16652
rect 18272 16612 18314 16652
rect 18354 16612 18396 16652
rect 18436 16612 18478 16652
rect 18518 16612 18560 16652
rect 18600 16612 33352 16652
rect 33392 16612 33434 16652
rect 33474 16612 33516 16652
rect 33556 16612 33598 16652
rect 33638 16612 33680 16652
rect 33720 16612 48472 16652
rect 48512 16612 48554 16652
rect 48594 16612 48636 16652
rect 48676 16612 48718 16652
rect 48758 16612 48800 16652
rect 48840 16612 63592 16652
rect 63632 16612 63674 16652
rect 63714 16612 63756 16652
rect 63796 16612 63838 16652
rect 63878 16612 63920 16652
rect 63960 16612 78712 16652
rect 78752 16612 78794 16652
rect 78834 16612 78876 16652
rect 78916 16612 78958 16652
rect 78998 16612 79040 16652
rect 79080 16612 93832 16652
rect 93872 16612 93914 16652
rect 93954 16612 93996 16652
rect 94036 16612 94078 16652
rect 94118 16612 94160 16652
rect 94200 16612 99360 16652
rect 576 16588 99360 16612
rect 651 16400 693 16409
rect 651 16360 652 16400
rect 692 16360 693 16400
rect 651 16351 693 16360
rect 33963 16400 34005 16409
rect 33963 16360 33964 16400
rect 34004 16360 34005 16400
rect 33963 16351 34005 16360
rect 33867 16316 33909 16325
rect 33867 16276 33868 16316
rect 33908 16276 33909 16316
rect 33867 16267 33909 16276
rect 34059 16316 34101 16325
rect 34059 16276 34060 16316
rect 34100 16276 34101 16316
rect 34059 16267 34101 16276
rect 33763 16232 33821 16233
rect 33763 16192 33772 16232
rect 33812 16192 33821 16232
rect 33763 16191 33821 16192
rect 34155 16232 34197 16241
rect 34155 16192 34156 16232
rect 34196 16192 34197 16232
rect 34155 16183 34197 16192
rect 37227 16232 37269 16241
rect 37227 16192 37228 16232
rect 37268 16192 37269 16232
rect 37227 16183 37269 16192
rect 37323 16232 37365 16241
rect 37323 16192 37324 16232
rect 37364 16192 37365 16232
rect 37323 16183 37365 16192
rect 38571 16232 38613 16241
rect 38571 16192 38572 16232
rect 38612 16192 38613 16232
rect 38571 16183 38613 16192
rect 39235 16232 39293 16233
rect 39235 16192 39244 16232
rect 39284 16192 39293 16232
rect 39235 16191 39293 16192
rect 37027 16064 37085 16065
rect 37027 16024 37036 16064
rect 37076 16024 37085 16064
rect 37027 16023 37085 16024
rect 576 15896 99360 15920
rect 576 15856 4352 15896
rect 4392 15856 4434 15896
rect 4474 15856 4516 15896
rect 4556 15856 4598 15896
rect 4638 15856 4680 15896
rect 4720 15856 19472 15896
rect 19512 15856 19554 15896
rect 19594 15856 19636 15896
rect 19676 15856 19718 15896
rect 19758 15856 19800 15896
rect 19840 15856 34592 15896
rect 34632 15856 34674 15896
rect 34714 15856 34756 15896
rect 34796 15856 34838 15896
rect 34878 15856 34920 15896
rect 34960 15856 49712 15896
rect 49752 15856 49794 15896
rect 49834 15856 49876 15896
rect 49916 15856 49958 15896
rect 49998 15856 50040 15896
rect 50080 15856 64832 15896
rect 64872 15856 64914 15896
rect 64954 15856 64996 15896
rect 65036 15856 65078 15896
rect 65118 15856 65160 15896
rect 65200 15856 79952 15896
rect 79992 15856 80034 15896
rect 80074 15856 80116 15896
rect 80156 15856 80198 15896
rect 80238 15856 80280 15896
rect 80320 15856 95072 15896
rect 95112 15856 95154 15896
rect 95194 15856 95236 15896
rect 95276 15856 95318 15896
rect 95358 15856 95400 15896
rect 95440 15856 99360 15896
rect 576 15832 99360 15856
rect 643 15728 701 15729
rect 643 15688 652 15728
rect 692 15688 701 15728
rect 643 15687 701 15688
rect 17827 15728 17885 15729
rect 17827 15688 17836 15728
rect 17876 15688 17885 15728
rect 17827 15687 17885 15688
rect 18211 15728 18269 15729
rect 18211 15688 18220 15728
rect 18260 15688 18269 15728
rect 18211 15687 18269 15688
rect 40003 15728 40061 15729
rect 40003 15688 40012 15728
rect 40052 15688 40061 15728
rect 40003 15687 40061 15688
rect 15435 15644 15477 15653
rect 15435 15604 15436 15644
rect 15476 15604 15477 15644
rect 15435 15595 15477 15604
rect 37611 15644 37653 15653
rect 37611 15604 37612 15644
rect 37652 15604 37653 15644
rect 37611 15595 37653 15604
rect 15811 15560 15869 15561
rect 15811 15520 15820 15560
rect 15860 15520 15869 15560
rect 15811 15519 15869 15520
rect 16675 15560 16733 15561
rect 16675 15520 16684 15560
rect 16724 15520 16733 15560
rect 16675 15519 16733 15520
rect 18307 15560 18365 15561
rect 18307 15520 18316 15560
rect 18356 15520 18365 15560
rect 18307 15519 18365 15520
rect 27907 15560 27965 15561
rect 27907 15520 27916 15560
rect 27956 15520 27965 15560
rect 27907 15519 27965 15520
rect 28299 15560 28341 15569
rect 28299 15520 28300 15560
rect 28340 15520 28341 15560
rect 28299 15511 28341 15520
rect 37987 15560 38045 15561
rect 37987 15520 37996 15560
rect 38036 15520 38045 15560
rect 37987 15519 38045 15520
rect 38851 15560 38909 15561
rect 38851 15520 38860 15560
rect 38900 15520 38909 15560
rect 38851 15519 38909 15520
rect 18883 15476 18941 15477
rect 18883 15436 18892 15476
rect 18932 15436 18941 15476
rect 18883 15435 18941 15436
rect 28011 15476 28053 15485
rect 28011 15436 28012 15476
rect 28052 15436 28053 15476
rect 28011 15427 28053 15436
rect 28203 15476 28245 15485
rect 28203 15436 28204 15476
rect 28244 15436 28245 15476
rect 28203 15427 28245 15436
rect 18499 15392 18557 15393
rect 18499 15352 18508 15392
rect 18548 15352 18557 15392
rect 18499 15351 18557 15352
rect 28107 15392 28149 15401
rect 28107 15352 28108 15392
rect 28148 15352 28149 15392
rect 28107 15343 28149 15352
rect 18699 15308 18741 15317
rect 18699 15268 18700 15308
rect 18740 15268 18741 15308
rect 18699 15259 18741 15268
rect 576 15140 99360 15164
rect 576 15100 3112 15140
rect 3152 15100 3194 15140
rect 3234 15100 3276 15140
rect 3316 15100 3358 15140
rect 3398 15100 3440 15140
rect 3480 15100 18232 15140
rect 18272 15100 18314 15140
rect 18354 15100 18396 15140
rect 18436 15100 18478 15140
rect 18518 15100 18560 15140
rect 18600 15100 33352 15140
rect 33392 15100 33434 15140
rect 33474 15100 33516 15140
rect 33556 15100 33598 15140
rect 33638 15100 33680 15140
rect 33720 15100 48472 15140
rect 48512 15100 48554 15140
rect 48594 15100 48636 15140
rect 48676 15100 48718 15140
rect 48758 15100 48800 15140
rect 48840 15100 63592 15140
rect 63632 15100 63674 15140
rect 63714 15100 63756 15140
rect 63796 15100 63838 15140
rect 63878 15100 63920 15140
rect 63960 15100 78712 15140
rect 78752 15100 78794 15140
rect 78834 15100 78876 15140
rect 78916 15100 78958 15140
rect 78998 15100 79040 15140
rect 79080 15100 93832 15140
rect 93872 15100 93914 15140
rect 93954 15100 93996 15140
rect 94036 15100 94078 15140
rect 94118 15100 94160 15140
rect 94200 15100 99360 15140
rect 576 15076 99360 15100
rect 25027 14972 25085 14973
rect 25027 14932 25036 14972
rect 25076 14932 25085 14972
rect 25027 14931 25085 14932
rect 22635 14720 22677 14729
rect 22635 14680 22636 14720
rect 22676 14680 22677 14720
rect 22635 14671 22677 14680
rect 23011 14720 23069 14721
rect 23011 14680 23020 14720
rect 23060 14680 23069 14720
rect 23011 14679 23069 14680
rect 23875 14720 23933 14721
rect 23875 14680 23884 14720
rect 23924 14680 23933 14720
rect 23875 14679 23933 14680
rect 643 14552 701 14553
rect 643 14512 652 14552
rect 692 14512 701 14552
rect 643 14511 701 14512
rect 576 14384 99360 14408
rect 576 14344 4352 14384
rect 4392 14344 4434 14384
rect 4474 14344 4516 14384
rect 4556 14344 4598 14384
rect 4638 14344 4680 14384
rect 4720 14344 19472 14384
rect 19512 14344 19554 14384
rect 19594 14344 19636 14384
rect 19676 14344 19718 14384
rect 19758 14344 19800 14384
rect 19840 14344 34592 14384
rect 34632 14344 34674 14384
rect 34714 14344 34756 14384
rect 34796 14344 34838 14384
rect 34878 14344 34920 14384
rect 34960 14344 49712 14384
rect 49752 14344 49794 14384
rect 49834 14344 49876 14384
rect 49916 14344 49958 14384
rect 49998 14344 50040 14384
rect 50080 14344 64832 14384
rect 64872 14344 64914 14384
rect 64954 14344 64996 14384
rect 65036 14344 65078 14384
rect 65118 14344 65160 14384
rect 65200 14344 79952 14384
rect 79992 14344 80034 14384
rect 80074 14344 80116 14384
rect 80156 14344 80198 14384
rect 80238 14344 80280 14384
rect 80320 14344 95072 14384
rect 95112 14344 95154 14384
rect 95194 14344 95236 14384
rect 95276 14344 95318 14384
rect 95358 14344 95400 14384
rect 95440 14344 99360 14384
rect 576 14320 99360 14344
rect 576 13628 99360 13652
rect 576 13588 3112 13628
rect 3152 13588 3194 13628
rect 3234 13588 3276 13628
rect 3316 13588 3358 13628
rect 3398 13588 3440 13628
rect 3480 13588 18232 13628
rect 18272 13588 18314 13628
rect 18354 13588 18396 13628
rect 18436 13588 18478 13628
rect 18518 13588 18560 13628
rect 18600 13588 33352 13628
rect 33392 13588 33434 13628
rect 33474 13588 33516 13628
rect 33556 13588 33598 13628
rect 33638 13588 33680 13628
rect 33720 13588 48472 13628
rect 48512 13588 48554 13628
rect 48594 13588 48636 13628
rect 48676 13588 48718 13628
rect 48758 13588 48800 13628
rect 48840 13588 63592 13628
rect 63632 13588 63674 13628
rect 63714 13588 63756 13628
rect 63796 13588 63838 13628
rect 63878 13588 63920 13628
rect 63960 13588 78712 13628
rect 78752 13588 78794 13628
rect 78834 13588 78876 13628
rect 78916 13588 78958 13628
rect 78998 13588 79040 13628
rect 79080 13588 93832 13628
rect 93872 13588 93914 13628
rect 93954 13588 93996 13628
rect 94036 13588 94078 13628
rect 94118 13588 94160 13628
rect 94200 13588 99360 13628
rect 576 13564 99360 13588
rect 33187 13208 33245 13209
rect 33187 13168 33196 13208
rect 33236 13168 33245 13208
rect 33187 13167 33245 13168
rect 643 13040 701 13041
rect 643 13000 652 13040
rect 692 13000 701 13040
rect 643 12999 701 13000
rect 32995 13040 33053 13041
rect 32995 13000 33004 13040
rect 33044 13000 33053 13040
rect 32995 12999 33053 13000
rect 33283 13040 33341 13041
rect 33283 13000 33292 13040
rect 33332 13000 33341 13040
rect 33283 12999 33341 13000
rect 576 12872 99360 12896
rect 576 12832 4352 12872
rect 4392 12832 4434 12872
rect 4474 12832 4516 12872
rect 4556 12832 4598 12872
rect 4638 12832 4680 12872
rect 4720 12832 19472 12872
rect 19512 12832 19554 12872
rect 19594 12832 19636 12872
rect 19676 12832 19718 12872
rect 19758 12832 19800 12872
rect 19840 12832 34592 12872
rect 34632 12832 34674 12872
rect 34714 12832 34756 12872
rect 34796 12832 34838 12872
rect 34878 12832 34920 12872
rect 34960 12832 49712 12872
rect 49752 12832 49794 12872
rect 49834 12832 49876 12872
rect 49916 12832 49958 12872
rect 49998 12832 50040 12872
rect 50080 12832 64832 12872
rect 64872 12832 64914 12872
rect 64954 12832 64996 12872
rect 65036 12832 65078 12872
rect 65118 12832 65160 12872
rect 65200 12832 79952 12872
rect 79992 12832 80034 12872
rect 80074 12832 80116 12872
rect 80156 12832 80198 12872
rect 80238 12832 80280 12872
rect 80320 12832 95072 12872
rect 95112 12832 95154 12872
rect 95194 12832 95236 12872
rect 95276 12832 95318 12872
rect 95358 12832 95400 12872
rect 95440 12832 99360 12872
rect 576 12808 99360 12832
rect 643 12704 701 12705
rect 643 12664 652 12704
rect 692 12664 701 12704
rect 643 12663 701 12664
rect 17739 12620 17781 12629
rect 17739 12580 17740 12620
rect 17780 12580 17781 12620
rect 17739 12571 17781 12580
rect 26475 12620 26517 12629
rect 26475 12580 26476 12620
rect 26516 12580 26517 12620
rect 26475 12571 26517 12580
rect 26859 12620 26901 12629
rect 26859 12580 26860 12620
rect 26900 12580 26901 12620
rect 26859 12571 26901 12580
rect 18115 12536 18173 12537
rect 18115 12496 18124 12536
rect 18164 12496 18173 12536
rect 18115 12495 18173 12496
rect 18979 12536 19037 12537
rect 18979 12496 18988 12536
rect 19028 12496 19037 12536
rect 18979 12495 19037 12496
rect 26371 12536 26429 12537
rect 26371 12496 26380 12536
rect 26420 12496 26429 12536
rect 26371 12495 26429 12496
rect 26571 12536 26613 12545
rect 26571 12496 26572 12536
rect 26612 12496 26613 12536
rect 26571 12487 26613 12496
rect 26755 12536 26813 12537
rect 26755 12496 26764 12536
rect 26804 12496 26813 12536
rect 26755 12495 26813 12496
rect 26955 12536 26997 12545
rect 26955 12496 26956 12536
rect 26996 12496 26997 12536
rect 26955 12487 26997 12496
rect 27243 12536 27285 12545
rect 27243 12496 27244 12536
rect 27284 12496 27285 12536
rect 27243 12487 27285 12496
rect 27819 12536 27861 12545
rect 27819 12496 27820 12536
rect 27860 12496 27861 12536
rect 27819 12487 27861 12496
rect 30891 12536 30933 12545
rect 30891 12496 30892 12536
rect 30932 12496 30933 12536
rect 30891 12487 30933 12496
rect 31267 12536 31325 12537
rect 31267 12496 31276 12536
rect 31316 12496 31325 12536
rect 31267 12495 31325 12496
rect 32131 12536 32189 12537
rect 32131 12496 32140 12536
rect 32180 12496 32189 12536
rect 32131 12495 32189 12496
rect 33291 12536 33333 12545
rect 33291 12496 33292 12536
rect 33332 12496 33333 12536
rect 33291 12487 33333 12496
rect 27435 12452 27477 12461
rect 27435 12412 27436 12452
rect 27476 12412 27477 12452
rect 27435 12403 27477 12412
rect 28011 12452 28053 12461
rect 28011 12412 28012 12452
rect 28052 12412 28053 12452
rect 28011 12403 28053 12412
rect 30699 12368 30741 12377
rect 30699 12328 30700 12368
rect 30740 12328 30741 12368
rect 30699 12319 30741 12328
rect 20131 12284 20189 12285
rect 20131 12244 20140 12284
rect 20180 12244 20189 12284
rect 20131 12243 20189 12244
rect 27243 12284 27285 12293
rect 27243 12244 27244 12284
rect 27284 12244 27285 12284
rect 27243 12235 27285 12244
rect 27819 12284 27861 12293
rect 27819 12244 27820 12284
rect 27860 12244 27861 12284
rect 27819 12235 27861 12244
rect 576 12116 99360 12140
rect 576 12076 3112 12116
rect 3152 12076 3194 12116
rect 3234 12076 3276 12116
rect 3316 12076 3358 12116
rect 3398 12076 3440 12116
rect 3480 12076 18232 12116
rect 18272 12076 18314 12116
rect 18354 12076 18396 12116
rect 18436 12076 18478 12116
rect 18518 12076 18560 12116
rect 18600 12076 33352 12116
rect 33392 12076 33434 12116
rect 33474 12076 33516 12116
rect 33556 12076 33598 12116
rect 33638 12076 33680 12116
rect 33720 12076 48472 12116
rect 48512 12076 48554 12116
rect 48594 12076 48636 12116
rect 48676 12076 48718 12116
rect 48758 12076 48800 12116
rect 48840 12076 63592 12116
rect 63632 12076 63674 12116
rect 63714 12076 63756 12116
rect 63796 12076 63838 12116
rect 63878 12076 63920 12116
rect 63960 12076 78712 12116
rect 78752 12076 78794 12116
rect 78834 12076 78876 12116
rect 78916 12076 78958 12116
rect 78998 12076 79040 12116
rect 79080 12076 93832 12116
rect 93872 12076 93914 12116
rect 93954 12076 93996 12116
rect 94036 12076 94078 12116
rect 94118 12076 94160 12116
rect 94200 12076 99360 12116
rect 576 12052 99360 12076
rect 24931 11948 24989 11949
rect 24931 11908 24940 11948
rect 24980 11908 24989 11948
rect 24931 11907 24989 11908
rect 835 11780 893 11781
rect 835 11740 844 11780
rect 884 11740 893 11780
rect 835 11739 893 11740
rect 22539 11696 22581 11705
rect 22539 11656 22540 11696
rect 22580 11656 22581 11696
rect 22539 11647 22581 11656
rect 22915 11696 22973 11697
rect 22915 11656 22924 11696
rect 22964 11656 22973 11696
rect 22915 11655 22973 11656
rect 23779 11696 23837 11697
rect 23779 11656 23788 11696
rect 23828 11656 23837 11696
rect 23779 11655 23837 11656
rect 651 11528 693 11537
rect 651 11488 652 11528
rect 692 11488 693 11528
rect 651 11479 693 11488
rect 576 11360 99360 11384
rect 576 11320 4352 11360
rect 4392 11320 4434 11360
rect 4474 11320 4516 11360
rect 4556 11320 4598 11360
rect 4638 11320 4680 11360
rect 4720 11320 19472 11360
rect 19512 11320 19554 11360
rect 19594 11320 19636 11360
rect 19676 11320 19718 11360
rect 19758 11320 19800 11360
rect 19840 11320 34592 11360
rect 34632 11320 34674 11360
rect 34714 11320 34756 11360
rect 34796 11320 34838 11360
rect 34878 11320 34920 11360
rect 34960 11320 49712 11360
rect 49752 11320 49794 11360
rect 49834 11320 49876 11360
rect 49916 11320 49958 11360
rect 49998 11320 50040 11360
rect 50080 11320 64832 11360
rect 64872 11320 64914 11360
rect 64954 11320 64996 11360
rect 65036 11320 65078 11360
rect 65118 11320 65160 11360
rect 65200 11320 79952 11360
rect 79992 11320 80034 11360
rect 80074 11320 80116 11360
rect 80156 11320 80198 11360
rect 80238 11320 80280 11360
rect 80320 11320 95072 11360
rect 95112 11320 95154 11360
rect 95194 11320 95236 11360
rect 95276 11320 95318 11360
rect 95358 11320 95400 11360
rect 95440 11320 99360 11360
rect 576 11296 99360 11320
rect 835 10940 893 10941
rect 835 10900 844 10940
rect 884 10900 893 10940
rect 835 10899 893 10900
rect 651 10772 693 10781
rect 651 10732 652 10772
rect 692 10732 693 10772
rect 651 10723 693 10732
rect 576 10604 99360 10628
rect 576 10564 3112 10604
rect 3152 10564 3194 10604
rect 3234 10564 3276 10604
rect 3316 10564 3358 10604
rect 3398 10564 3440 10604
rect 3480 10564 18232 10604
rect 18272 10564 18314 10604
rect 18354 10564 18396 10604
rect 18436 10564 18478 10604
rect 18518 10564 18560 10604
rect 18600 10564 33352 10604
rect 33392 10564 33434 10604
rect 33474 10564 33516 10604
rect 33556 10564 33598 10604
rect 33638 10564 33680 10604
rect 33720 10564 48472 10604
rect 48512 10564 48554 10604
rect 48594 10564 48636 10604
rect 48676 10564 48718 10604
rect 48758 10564 48800 10604
rect 48840 10564 63592 10604
rect 63632 10564 63674 10604
rect 63714 10564 63756 10604
rect 63796 10564 63838 10604
rect 63878 10564 63920 10604
rect 63960 10564 78712 10604
rect 78752 10564 78794 10604
rect 78834 10564 78876 10604
rect 78916 10564 78958 10604
rect 78998 10564 79040 10604
rect 79080 10564 93832 10604
rect 93872 10564 93914 10604
rect 93954 10564 93996 10604
rect 94036 10564 94078 10604
rect 94118 10564 94160 10604
rect 94200 10564 99360 10604
rect 576 10540 99360 10564
rect 835 10268 893 10269
rect 835 10228 844 10268
rect 884 10228 893 10268
rect 835 10227 893 10228
rect 651 10016 693 10025
rect 651 9976 652 10016
rect 692 9976 693 10016
rect 651 9967 693 9976
rect 576 9848 99360 9872
rect 576 9808 4352 9848
rect 4392 9808 4434 9848
rect 4474 9808 4516 9848
rect 4556 9808 4598 9848
rect 4638 9808 4680 9848
rect 4720 9808 19472 9848
rect 19512 9808 19554 9848
rect 19594 9808 19636 9848
rect 19676 9808 19718 9848
rect 19758 9808 19800 9848
rect 19840 9808 34592 9848
rect 34632 9808 34674 9848
rect 34714 9808 34756 9848
rect 34796 9808 34838 9848
rect 34878 9808 34920 9848
rect 34960 9808 49712 9848
rect 49752 9808 49794 9848
rect 49834 9808 49876 9848
rect 49916 9808 49958 9848
rect 49998 9808 50040 9848
rect 50080 9808 64832 9848
rect 64872 9808 64914 9848
rect 64954 9808 64996 9848
rect 65036 9808 65078 9848
rect 65118 9808 65160 9848
rect 65200 9808 79952 9848
rect 79992 9808 80034 9848
rect 80074 9808 80116 9848
rect 80156 9808 80198 9848
rect 80238 9808 80280 9848
rect 80320 9808 95072 9848
rect 95112 9808 95154 9848
rect 95194 9808 95236 9848
rect 95276 9808 95318 9848
rect 95358 9808 95400 9848
rect 95440 9808 99360 9848
rect 576 9784 99360 9808
rect 835 9428 893 9429
rect 835 9388 844 9428
rect 884 9388 893 9428
rect 835 9387 893 9388
rect 651 9260 693 9269
rect 651 9220 652 9260
rect 692 9220 693 9260
rect 651 9211 693 9220
rect 576 9092 99360 9116
rect 576 9052 3112 9092
rect 3152 9052 3194 9092
rect 3234 9052 3276 9092
rect 3316 9052 3358 9092
rect 3398 9052 3440 9092
rect 3480 9052 18232 9092
rect 18272 9052 18314 9092
rect 18354 9052 18396 9092
rect 18436 9052 18478 9092
rect 18518 9052 18560 9092
rect 18600 9052 33352 9092
rect 33392 9052 33434 9092
rect 33474 9052 33516 9092
rect 33556 9052 33598 9092
rect 33638 9052 33680 9092
rect 33720 9052 48472 9092
rect 48512 9052 48554 9092
rect 48594 9052 48636 9092
rect 48676 9052 48718 9092
rect 48758 9052 48800 9092
rect 48840 9052 63592 9092
rect 63632 9052 63674 9092
rect 63714 9052 63756 9092
rect 63796 9052 63838 9092
rect 63878 9052 63920 9092
rect 63960 9052 78712 9092
rect 78752 9052 78794 9092
rect 78834 9052 78876 9092
rect 78916 9052 78958 9092
rect 78998 9052 79040 9092
rect 79080 9052 93832 9092
rect 93872 9052 93914 9092
rect 93954 9052 93996 9092
rect 94036 9052 94078 9092
rect 94118 9052 94160 9092
rect 94200 9052 99360 9092
rect 576 9028 99360 9052
rect 835 8756 893 8757
rect 835 8716 844 8756
rect 884 8716 893 8756
rect 835 8715 893 8716
rect 651 8504 693 8513
rect 651 8464 652 8504
rect 692 8464 693 8504
rect 651 8455 693 8464
rect 576 8336 99360 8360
rect 576 8296 4352 8336
rect 4392 8296 4434 8336
rect 4474 8296 4516 8336
rect 4556 8296 4598 8336
rect 4638 8296 4680 8336
rect 4720 8296 19472 8336
rect 19512 8296 19554 8336
rect 19594 8296 19636 8336
rect 19676 8296 19718 8336
rect 19758 8296 19800 8336
rect 19840 8296 34592 8336
rect 34632 8296 34674 8336
rect 34714 8296 34756 8336
rect 34796 8296 34838 8336
rect 34878 8296 34920 8336
rect 34960 8296 49712 8336
rect 49752 8296 49794 8336
rect 49834 8296 49876 8336
rect 49916 8296 49958 8336
rect 49998 8296 50040 8336
rect 50080 8296 64832 8336
rect 64872 8296 64914 8336
rect 64954 8296 64996 8336
rect 65036 8296 65078 8336
rect 65118 8296 65160 8336
rect 65200 8296 79952 8336
rect 79992 8296 80034 8336
rect 80074 8296 80116 8336
rect 80156 8296 80198 8336
rect 80238 8296 80280 8336
rect 80320 8296 95072 8336
rect 95112 8296 95154 8336
rect 95194 8296 95236 8336
rect 95276 8296 95318 8336
rect 95358 8296 95400 8336
rect 95440 8296 99360 8336
rect 576 8272 99360 8296
rect 835 7916 893 7917
rect 835 7876 844 7916
rect 884 7876 893 7916
rect 835 7875 893 7876
rect 651 7748 693 7757
rect 651 7708 652 7748
rect 692 7708 693 7748
rect 651 7699 693 7708
rect 576 7580 99360 7604
rect 576 7540 3112 7580
rect 3152 7540 3194 7580
rect 3234 7540 3276 7580
rect 3316 7540 3358 7580
rect 3398 7540 3440 7580
rect 3480 7540 18232 7580
rect 18272 7540 18314 7580
rect 18354 7540 18396 7580
rect 18436 7540 18478 7580
rect 18518 7540 18560 7580
rect 18600 7540 33352 7580
rect 33392 7540 33434 7580
rect 33474 7540 33516 7580
rect 33556 7540 33598 7580
rect 33638 7540 33680 7580
rect 33720 7540 48472 7580
rect 48512 7540 48554 7580
rect 48594 7540 48636 7580
rect 48676 7540 48718 7580
rect 48758 7540 48800 7580
rect 48840 7540 63592 7580
rect 63632 7540 63674 7580
rect 63714 7540 63756 7580
rect 63796 7540 63838 7580
rect 63878 7540 63920 7580
rect 63960 7540 78712 7580
rect 78752 7540 78794 7580
rect 78834 7540 78876 7580
rect 78916 7540 78958 7580
rect 78998 7540 79040 7580
rect 79080 7540 93832 7580
rect 93872 7540 93914 7580
rect 93954 7540 93996 7580
rect 94036 7540 94078 7580
rect 94118 7540 94160 7580
rect 94200 7540 99360 7580
rect 576 7516 99360 7540
rect 835 7244 893 7245
rect 835 7204 844 7244
rect 884 7204 893 7244
rect 835 7203 893 7204
rect 651 6992 693 7001
rect 651 6952 652 6992
rect 692 6952 693 6992
rect 651 6943 693 6952
rect 576 6824 99360 6848
rect 576 6784 4352 6824
rect 4392 6784 4434 6824
rect 4474 6784 4516 6824
rect 4556 6784 4598 6824
rect 4638 6784 4680 6824
rect 4720 6784 19472 6824
rect 19512 6784 19554 6824
rect 19594 6784 19636 6824
rect 19676 6784 19718 6824
rect 19758 6784 19800 6824
rect 19840 6784 34592 6824
rect 34632 6784 34674 6824
rect 34714 6784 34756 6824
rect 34796 6784 34838 6824
rect 34878 6784 34920 6824
rect 34960 6784 49712 6824
rect 49752 6784 49794 6824
rect 49834 6784 49876 6824
rect 49916 6784 49958 6824
rect 49998 6784 50040 6824
rect 50080 6784 64832 6824
rect 64872 6784 64914 6824
rect 64954 6784 64996 6824
rect 65036 6784 65078 6824
rect 65118 6784 65160 6824
rect 65200 6784 79952 6824
rect 79992 6784 80034 6824
rect 80074 6784 80116 6824
rect 80156 6784 80198 6824
rect 80238 6784 80280 6824
rect 80320 6784 95072 6824
rect 95112 6784 95154 6824
rect 95194 6784 95236 6824
rect 95276 6784 95318 6824
rect 95358 6784 95400 6824
rect 95440 6784 99360 6824
rect 576 6760 99360 6784
rect 576 6068 99360 6092
rect 576 6028 3112 6068
rect 3152 6028 3194 6068
rect 3234 6028 3276 6068
rect 3316 6028 3358 6068
rect 3398 6028 3440 6068
rect 3480 6028 18232 6068
rect 18272 6028 18314 6068
rect 18354 6028 18396 6068
rect 18436 6028 18478 6068
rect 18518 6028 18560 6068
rect 18600 6028 33352 6068
rect 33392 6028 33434 6068
rect 33474 6028 33516 6068
rect 33556 6028 33598 6068
rect 33638 6028 33680 6068
rect 33720 6028 48472 6068
rect 48512 6028 48554 6068
rect 48594 6028 48636 6068
rect 48676 6028 48718 6068
rect 48758 6028 48800 6068
rect 48840 6028 63592 6068
rect 63632 6028 63674 6068
rect 63714 6028 63756 6068
rect 63796 6028 63838 6068
rect 63878 6028 63920 6068
rect 63960 6028 78712 6068
rect 78752 6028 78794 6068
rect 78834 6028 78876 6068
rect 78916 6028 78958 6068
rect 78998 6028 79040 6068
rect 79080 6028 93832 6068
rect 93872 6028 93914 6068
rect 93954 6028 93996 6068
rect 94036 6028 94078 6068
rect 94118 6028 94160 6068
rect 94200 6028 99360 6068
rect 576 6004 99360 6028
rect 835 5732 893 5733
rect 835 5692 844 5732
rect 884 5692 893 5732
rect 835 5691 893 5692
rect 651 5480 693 5489
rect 651 5440 652 5480
rect 692 5440 693 5480
rect 651 5431 693 5440
rect 576 5312 99360 5336
rect 576 5272 4352 5312
rect 4392 5272 4434 5312
rect 4474 5272 4516 5312
rect 4556 5272 4598 5312
rect 4638 5272 4680 5312
rect 4720 5272 19472 5312
rect 19512 5272 19554 5312
rect 19594 5272 19636 5312
rect 19676 5272 19718 5312
rect 19758 5272 19800 5312
rect 19840 5272 34592 5312
rect 34632 5272 34674 5312
rect 34714 5272 34756 5312
rect 34796 5272 34838 5312
rect 34878 5272 34920 5312
rect 34960 5272 49712 5312
rect 49752 5272 49794 5312
rect 49834 5272 49876 5312
rect 49916 5272 49958 5312
rect 49998 5272 50040 5312
rect 50080 5272 64832 5312
rect 64872 5272 64914 5312
rect 64954 5272 64996 5312
rect 65036 5272 65078 5312
rect 65118 5272 65160 5312
rect 65200 5272 79952 5312
rect 79992 5272 80034 5312
rect 80074 5272 80116 5312
rect 80156 5272 80198 5312
rect 80238 5272 80280 5312
rect 80320 5272 95072 5312
rect 95112 5272 95154 5312
rect 95194 5272 95236 5312
rect 95276 5272 95318 5312
rect 95358 5272 95400 5312
rect 95440 5272 99360 5312
rect 576 5248 99360 5272
rect 835 4892 893 4893
rect 835 4852 844 4892
rect 884 4852 893 4892
rect 835 4851 893 4852
rect 651 4808 693 4817
rect 651 4768 652 4808
rect 692 4768 693 4808
rect 651 4759 693 4768
rect 576 4556 99360 4580
rect 576 4516 3112 4556
rect 3152 4516 3194 4556
rect 3234 4516 3276 4556
rect 3316 4516 3358 4556
rect 3398 4516 3440 4556
rect 3480 4516 18232 4556
rect 18272 4516 18314 4556
rect 18354 4516 18396 4556
rect 18436 4516 18478 4556
rect 18518 4516 18560 4556
rect 18600 4516 33352 4556
rect 33392 4516 33434 4556
rect 33474 4516 33516 4556
rect 33556 4516 33598 4556
rect 33638 4516 33680 4556
rect 33720 4516 48472 4556
rect 48512 4516 48554 4556
rect 48594 4516 48636 4556
rect 48676 4516 48718 4556
rect 48758 4516 48800 4556
rect 48840 4516 63592 4556
rect 63632 4516 63674 4556
rect 63714 4516 63756 4556
rect 63796 4516 63838 4556
rect 63878 4516 63920 4556
rect 63960 4516 78712 4556
rect 78752 4516 78794 4556
rect 78834 4516 78876 4556
rect 78916 4516 78958 4556
rect 78998 4516 79040 4556
rect 79080 4516 93832 4556
rect 93872 4516 93914 4556
rect 93954 4516 93996 4556
rect 94036 4516 94078 4556
rect 94118 4516 94160 4556
rect 94200 4516 99360 4556
rect 576 4492 99360 4516
rect 835 4220 893 4221
rect 835 4180 844 4220
rect 884 4180 893 4220
rect 835 4179 893 4180
rect 651 3968 693 3977
rect 651 3928 652 3968
rect 692 3928 693 3968
rect 651 3919 693 3928
rect 576 3800 99360 3824
rect 576 3760 4352 3800
rect 4392 3760 4434 3800
rect 4474 3760 4516 3800
rect 4556 3760 4598 3800
rect 4638 3760 4680 3800
rect 4720 3760 19472 3800
rect 19512 3760 19554 3800
rect 19594 3760 19636 3800
rect 19676 3760 19718 3800
rect 19758 3760 19800 3800
rect 19840 3760 34592 3800
rect 34632 3760 34674 3800
rect 34714 3760 34756 3800
rect 34796 3760 34838 3800
rect 34878 3760 34920 3800
rect 34960 3760 49712 3800
rect 49752 3760 49794 3800
rect 49834 3760 49876 3800
rect 49916 3760 49958 3800
rect 49998 3760 50040 3800
rect 50080 3760 64832 3800
rect 64872 3760 64914 3800
rect 64954 3760 64996 3800
rect 65036 3760 65078 3800
rect 65118 3760 65160 3800
rect 65200 3760 79952 3800
rect 79992 3760 80034 3800
rect 80074 3760 80116 3800
rect 80156 3760 80198 3800
rect 80238 3760 80280 3800
rect 80320 3760 95072 3800
rect 95112 3760 95154 3800
rect 95194 3760 95236 3800
rect 95276 3760 95318 3800
rect 95358 3760 95400 3800
rect 95440 3760 99360 3800
rect 576 3736 99360 3760
rect 835 3380 893 3381
rect 835 3340 844 3380
rect 884 3340 893 3380
rect 835 3339 893 3340
rect 651 3212 693 3221
rect 651 3172 652 3212
rect 692 3172 693 3212
rect 651 3163 693 3172
rect 576 3044 99360 3068
rect 576 3004 3112 3044
rect 3152 3004 3194 3044
rect 3234 3004 3276 3044
rect 3316 3004 3358 3044
rect 3398 3004 3440 3044
rect 3480 3004 18232 3044
rect 18272 3004 18314 3044
rect 18354 3004 18396 3044
rect 18436 3004 18478 3044
rect 18518 3004 18560 3044
rect 18600 3004 33352 3044
rect 33392 3004 33434 3044
rect 33474 3004 33516 3044
rect 33556 3004 33598 3044
rect 33638 3004 33680 3044
rect 33720 3004 48472 3044
rect 48512 3004 48554 3044
rect 48594 3004 48636 3044
rect 48676 3004 48718 3044
rect 48758 3004 48800 3044
rect 48840 3004 63592 3044
rect 63632 3004 63674 3044
rect 63714 3004 63756 3044
rect 63796 3004 63838 3044
rect 63878 3004 63920 3044
rect 63960 3004 78712 3044
rect 78752 3004 78794 3044
rect 78834 3004 78876 3044
rect 78916 3004 78958 3044
rect 78998 3004 79040 3044
rect 79080 3004 93832 3044
rect 93872 3004 93914 3044
rect 93954 3004 93996 3044
rect 94036 3004 94078 3044
rect 94118 3004 94160 3044
rect 94200 3004 99360 3044
rect 576 2980 99360 3004
rect 835 2708 893 2709
rect 835 2668 844 2708
rect 884 2668 893 2708
rect 835 2667 893 2668
rect 651 2456 693 2465
rect 651 2416 652 2456
rect 692 2416 693 2456
rect 651 2407 693 2416
rect 576 2288 99360 2312
rect 576 2248 4352 2288
rect 4392 2248 4434 2288
rect 4474 2248 4516 2288
rect 4556 2248 4598 2288
rect 4638 2248 4680 2288
rect 4720 2248 19472 2288
rect 19512 2248 19554 2288
rect 19594 2248 19636 2288
rect 19676 2248 19718 2288
rect 19758 2248 19800 2288
rect 19840 2248 34592 2288
rect 34632 2248 34674 2288
rect 34714 2248 34756 2288
rect 34796 2248 34838 2288
rect 34878 2248 34920 2288
rect 34960 2248 49712 2288
rect 49752 2248 49794 2288
rect 49834 2248 49876 2288
rect 49916 2248 49958 2288
rect 49998 2248 50040 2288
rect 50080 2248 64832 2288
rect 64872 2248 64914 2288
rect 64954 2248 64996 2288
rect 65036 2248 65078 2288
rect 65118 2248 65160 2288
rect 65200 2248 79952 2288
rect 79992 2248 80034 2288
rect 80074 2248 80116 2288
rect 80156 2248 80198 2288
rect 80238 2248 80280 2288
rect 80320 2248 95072 2288
rect 95112 2248 95154 2288
rect 95194 2248 95236 2288
rect 95276 2248 95318 2288
rect 95358 2248 95400 2288
rect 95440 2248 99360 2288
rect 576 2224 99360 2248
rect 576 1532 99360 1556
rect 576 1492 3112 1532
rect 3152 1492 3194 1532
rect 3234 1492 3276 1532
rect 3316 1492 3358 1532
rect 3398 1492 3440 1532
rect 3480 1492 18232 1532
rect 18272 1492 18314 1532
rect 18354 1492 18396 1532
rect 18436 1492 18478 1532
rect 18518 1492 18560 1532
rect 18600 1492 33352 1532
rect 33392 1492 33434 1532
rect 33474 1492 33516 1532
rect 33556 1492 33598 1532
rect 33638 1492 33680 1532
rect 33720 1492 48472 1532
rect 48512 1492 48554 1532
rect 48594 1492 48636 1532
rect 48676 1492 48718 1532
rect 48758 1492 48800 1532
rect 48840 1492 63592 1532
rect 63632 1492 63674 1532
rect 63714 1492 63756 1532
rect 63796 1492 63838 1532
rect 63878 1492 63920 1532
rect 63960 1492 78712 1532
rect 78752 1492 78794 1532
rect 78834 1492 78876 1532
rect 78916 1492 78958 1532
rect 78998 1492 79040 1532
rect 79080 1492 93832 1532
rect 93872 1492 93914 1532
rect 93954 1492 93996 1532
rect 94036 1492 94078 1532
rect 94118 1492 94160 1532
rect 94200 1492 99360 1532
rect 576 1468 99360 1492
rect 576 776 99360 800
rect 576 736 4352 776
rect 4392 736 4434 776
rect 4474 736 4516 776
rect 4556 736 4598 776
rect 4638 736 4680 776
rect 4720 736 19472 776
rect 19512 736 19554 776
rect 19594 736 19636 776
rect 19676 736 19718 776
rect 19758 736 19800 776
rect 19840 736 34592 776
rect 34632 736 34674 776
rect 34714 736 34756 776
rect 34796 736 34838 776
rect 34878 736 34920 776
rect 34960 736 49712 776
rect 49752 736 49794 776
rect 49834 736 49876 776
rect 49916 736 49958 776
rect 49998 736 50040 776
rect 50080 736 64832 776
rect 64872 736 64914 776
rect 64954 736 64996 776
rect 65036 736 65078 776
rect 65118 736 65160 776
rect 65200 736 79952 776
rect 79992 736 80034 776
rect 80074 736 80116 776
rect 80156 736 80198 776
rect 80238 736 80280 776
rect 80320 736 95072 776
rect 95112 736 95154 776
rect 95194 736 95236 776
rect 95276 736 95318 776
rect 95358 736 95400 776
rect 95440 736 99360 776
rect 576 712 99360 736
<< via1 >>
rect 4352 38536 4392 38576
rect 4434 38536 4474 38576
rect 4516 38536 4556 38576
rect 4598 38536 4638 38576
rect 4680 38536 4720 38576
rect 19472 38536 19512 38576
rect 19554 38536 19594 38576
rect 19636 38536 19676 38576
rect 19718 38536 19758 38576
rect 19800 38536 19840 38576
rect 34592 38536 34632 38576
rect 34674 38536 34714 38576
rect 34756 38536 34796 38576
rect 34838 38536 34878 38576
rect 34920 38536 34960 38576
rect 49712 38536 49752 38576
rect 49794 38536 49834 38576
rect 49876 38536 49916 38576
rect 49958 38536 49998 38576
rect 50040 38536 50080 38576
rect 64832 38536 64872 38576
rect 64914 38536 64954 38576
rect 64996 38536 65036 38576
rect 65078 38536 65118 38576
rect 65160 38536 65200 38576
rect 79952 38536 79992 38576
rect 80034 38536 80074 38576
rect 80116 38536 80156 38576
rect 80198 38536 80238 38576
rect 80280 38536 80320 38576
rect 95072 38536 95112 38576
rect 95154 38536 95194 38576
rect 95236 38536 95276 38576
rect 95318 38536 95358 38576
rect 95400 38536 95440 38576
rect 3112 37780 3152 37820
rect 3194 37780 3234 37820
rect 3276 37780 3316 37820
rect 3358 37780 3398 37820
rect 3440 37780 3480 37820
rect 18232 37780 18272 37820
rect 18314 37780 18354 37820
rect 18396 37780 18436 37820
rect 18478 37780 18518 37820
rect 18560 37780 18600 37820
rect 33352 37780 33392 37820
rect 33434 37780 33474 37820
rect 33516 37780 33556 37820
rect 33598 37780 33638 37820
rect 33680 37780 33720 37820
rect 48472 37780 48512 37820
rect 48554 37780 48594 37820
rect 48636 37780 48676 37820
rect 48718 37780 48758 37820
rect 48800 37780 48840 37820
rect 63592 37780 63632 37820
rect 63674 37780 63714 37820
rect 63756 37780 63796 37820
rect 63838 37780 63878 37820
rect 63920 37780 63960 37820
rect 78712 37780 78752 37820
rect 78794 37780 78834 37820
rect 78876 37780 78916 37820
rect 78958 37780 78998 37820
rect 79040 37780 79080 37820
rect 93832 37780 93872 37820
rect 93914 37780 93954 37820
rect 93996 37780 94036 37820
rect 94078 37780 94118 37820
rect 94160 37780 94200 37820
rect 4352 37024 4392 37064
rect 4434 37024 4474 37064
rect 4516 37024 4556 37064
rect 4598 37024 4638 37064
rect 4680 37024 4720 37064
rect 19472 37024 19512 37064
rect 19554 37024 19594 37064
rect 19636 37024 19676 37064
rect 19718 37024 19758 37064
rect 19800 37024 19840 37064
rect 34592 37024 34632 37064
rect 34674 37024 34714 37064
rect 34756 37024 34796 37064
rect 34838 37024 34878 37064
rect 34920 37024 34960 37064
rect 49712 37024 49752 37064
rect 49794 37024 49834 37064
rect 49876 37024 49916 37064
rect 49958 37024 49998 37064
rect 50040 37024 50080 37064
rect 64832 37024 64872 37064
rect 64914 37024 64954 37064
rect 64996 37024 65036 37064
rect 65078 37024 65118 37064
rect 65160 37024 65200 37064
rect 79952 37024 79992 37064
rect 80034 37024 80074 37064
rect 80116 37024 80156 37064
rect 80198 37024 80238 37064
rect 80280 37024 80320 37064
rect 95072 37024 95112 37064
rect 95154 37024 95194 37064
rect 95236 37024 95276 37064
rect 95318 37024 95358 37064
rect 95400 37024 95440 37064
rect 3112 36268 3152 36308
rect 3194 36268 3234 36308
rect 3276 36268 3316 36308
rect 3358 36268 3398 36308
rect 3440 36268 3480 36308
rect 18232 36268 18272 36308
rect 18314 36268 18354 36308
rect 18396 36268 18436 36308
rect 18478 36268 18518 36308
rect 18560 36268 18600 36308
rect 33352 36268 33392 36308
rect 33434 36268 33474 36308
rect 33516 36268 33556 36308
rect 33598 36268 33638 36308
rect 33680 36268 33720 36308
rect 48472 36268 48512 36308
rect 48554 36268 48594 36308
rect 48636 36268 48676 36308
rect 48718 36268 48758 36308
rect 48800 36268 48840 36308
rect 63592 36268 63632 36308
rect 63674 36268 63714 36308
rect 63756 36268 63796 36308
rect 63838 36268 63878 36308
rect 63920 36268 63960 36308
rect 78712 36268 78752 36308
rect 78794 36268 78834 36308
rect 78876 36268 78916 36308
rect 78958 36268 78998 36308
rect 79040 36268 79080 36308
rect 93832 36268 93872 36308
rect 93914 36268 93954 36308
rect 93996 36268 94036 36308
rect 94078 36268 94118 36308
rect 94160 36268 94200 36308
rect 4352 35512 4392 35552
rect 4434 35512 4474 35552
rect 4516 35512 4556 35552
rect 4598 35512 4638 35552
rect 4680 35512 4720 35552
rect 19472 35512 19512 35552
rect 19554 35512 19594 35552
rect 19636 35512 19676 35552
rect 19718 35512 19758 35552
rect 19800 35512 19840 35552
rect 34592 35512 34632 35552
rect 34674 35512 34714 35552
rect 34756 35512 34796 35552
rect 34838 35512 34878 35552
rect 34920 35512 34960 35552
rect 49712 35512 49752 35552
rect 49794 35512 49834 35552
rect 49876 35512 49916 35552
rect 49958 35512 49998 35552
rect 50040 35512 50080 35552
rect 64832 35512 64872 35552
rect 64914 35512 64954 35552
rect 64996 35512 65036 35552
rect 65078 35512 65118 35552
rect 65160 35512 65200 35552
rect 79952 35512 79992 35552
rect 80034 35512 80074 35552
rect 80116 35512 80156 35552
rect 80198 35512 80238 35552
rect 80280 35512 80320 35552
rect 95072 35512 95112 35552
rect 95154 35512 95194 35552
rect 95236 35512 95276 35552
rect 95318 35512 95358 35552
rect 95400 35512 95440 35552
rect 652 35176 692 35216
rect 844 35176 884 35216
rect 3112 34756 3152 34796
rect 3194 34756 3234 34796
rect 3276 34756 3316 34796
rect 3358 34756 3398 34796
rect 3440 34756 3480 34796
rect 18232 34756 18272 34796
rect 18314 34756 18354 34796
rect 18396 34756 18436 34796
rect 18478 34756 18518 34796
rect 18560 34756 18600 34796
rect 33352 34756 33392 34796
rect 33434 34756 33474 34796
rect 33516 34756 33556 34796
rect 33598 34756 33638 34796
rect 33680 34756 33720 34796
rect 48472 34756 48512 34796
rect 48554 34756 48594 34796
rect 48636 34756 48676 34796
rect 48718 34756 48758 34796
rect 48800 34756 48840 34796
rect 63592 34756 63632 34796
rect 63674 34756 63714 34796
rect 63756 34756 63796 34796
rect 63838 34756 63878 34796
rect 63920 34756 63960 34796
rect 78712 34756 78752 34796
rect 78794 34756 78834 34796
rect 78876 34756 78916 34796
rect 78958 34756 78998 34796
rect 79040 34756 79080 34796
rect 93832 34756 93872 34796
rect 93914 34756 93954 34796
rect 93996 34756 94036 34796
rect 94078 34756 94118 34796
rect 94160 34756 94200 34796
rect 652 34336 692 34376
rect 844 34336 884 34376
rect 4352 34000 4392 34040
rect 4434 34000 4474 34040
rect 4516 34000 4556 34040
rect 4598 34000 4638 34040
rect 4680 34000 4720 34040
rect 19472 34000 19512 34040
rect 19554 34000 19594 34040
rect 19636 34000 19676 34040
rect 19718 34000 19758 34040
rect 19800 34000 19840 34040
rect 34592 34000 34632 34040
rect 34674 34000 34714 34040
rect 34756 34000 34796 34040
rect 34838 34000 34878 34040
rect 34920 34000 34960 34040
rect 49712 34000 49752 34040
rect 49794 34000 49834 34040
rect 49876 34000 49916 34040
rect 49958 34000 49998 34040
rect 50040 34000 50080 34040
rect 64832 34000 64872 34040
rect 64914 34000 64954 34040
rect 64996 34000 65036 34040
rect 65078 34000 65118 34040
rect 65160 34000 65200 34040
rect 79952 34000 79992 34040
rect 80034 34000 80074 34040
rect 80116 34000 80156 34040
rect 80198 34000 80238 34040
rect 80280 34000 80320 34040
rect 95072 34000 95112 34040
rect 95154 34000 95194 34040
rect 95236 34000 95276 34040
rect 95318 34000 95358 34040
rect 95400 34000 95440 34040
rect 652 33664 692 33704
rect 844 33664 884 33704
rect 3112 33244 3152 33284
rect 3194 33244 3234 33284
rect 3276 33244 3316 33284
rect 3358 33244 3398 33284
rect 3440 33244 3480 33284
rect 18232 33244 18272 33284
rect 18314 33244 18354 33284
rect 18396 33244 18436 33284
rect 18478 33244 18518 33284
rect 18560 33244 18600 33284
rect 33352 33244 33392 33284
rect 33434 33244 33474 33284
rect 33516 33244 33556 33284
rect 33598 33244 33638 33284
rect 33680 33244 33720 33284
rect 48472 33244 48512 33284
rect 48554 33244 48594 33284
rect 48636 33244 48676 33284
rect 48718 33244 48758 33284
rect 48800 33244 48840 33284
rect 63592 33244 63632 33284
rect 63674 33244 63714 33284
rect 63756 33244 63796 33284
rect 63838 33244 63878 33284
rect 63920 33244 63960 33284
rect 78712 33244 78752 33284
rect 78794 33244 78834 33284
rect 78876 33244 78916 33284
rect 78958 33244 78998 33284
rect 79040 33244 79080 33284
rect 93832 33244 93872 33284
rect 93914 33244 93954 33284
rect 93996 33244 94036 33284
rect 94078 33244 94118 33284
rect 94160 33244 94200 33284
rect 652 32824 692 32864
rect 844 32824 884 32864
rect 4352 32488 4392 32528
rect 4434 32488 4474 32528
rect 4516 32488 4556 32528
rect 4598 32488 4638 32528
rect 4680 32488 4720 32528
rect 19472 32488 19512 32528
rect 19554 32488 19594 32528
rect 19636 32488 19676 32528
rect 19718 32488 19758 32528
rect 19800 32488 19840 32528
rect 34592 32488 34632 32528
rect 34674 32488 34714 32528
rect 34756 32488 34796 32528
rect 34838 32488 34878 32528
rect 34920 32488 34960 32528
rect 49712 32488 49752 32528
rect 49794 32488 49834 32528
rect 49876 32488 49916 32528
rect 49958 32488 49998 32528
rect 50040 32488 50080 32528
rect 64832 32488 64872 32528
rect 64914 32488 64954 32528
rect 64996 32488 65036 32528
rect 65078 32488 65118 32528
rect 65160 32488 65200 32528
rect 79952 32488 79992 32528
rect 80034 32488 80074 32528
rect 80116 32488 80156 32528
rect 80198 32488 80238 32528
rect 80280 32488 80320 32528
rect 95072 32488 95112 32528
rect 95154 32488 95194 32528
rect 95236 32488 95276 32528
rect 95318 32488 95358 32528
rect 95400 32488 95440 32528
rect 27436 32152 27476 32192
rect 652 32068 692 32108
rect 844 31900 884 31940
rect 27532 31900 27572 31940
rect 3112 31732 3152 31772
rect 3194 31732 3234 31772
rect 3276 31732 3316 31772
rect 3358 31732 3398 31772
rect 3440 31732 3480 31772
rect 18232 31732 18272 31772
rect 18314 31732 18354 31772
rect 18396 31732 18436 31772
rect 18478 31732 18518 31772
rect 18560 31732 18600 31772
rect 33352 31732 33392 31772
rect 33434 31732 33474 31772
rect 33516 31732 33556 31772
rect 33598 31732 33638 31772
rect 33680 31732 33720 31772
rect 48472 31732 48512 31772
rect 48554 31732 48594 31772
rect 48636 31732 48676 31772
rect 48718 31732 48758 31772
rect 48800 31732 48840 31772
rect 63592 31732 63632 31772
rect 63674 31732 63714 31772
rect 63756 31732 63796 31772
rect 63838 31732 63878 31772
rect 63920 31732 63960 31772
rect 78712 31732 78752 31772
rect 78794 31732 78834 31772
rect 78876 31732 78916 31772
rect 78958 31732 78998 31772
rect 79040 31732 79080 31772
rect 93832 31732 93872 31772
rect 93914 31732 93954 31772
rect 93996 31732 94036 31772
rect 94078 31732 94118 31772
rect 94160 31732 94200 31772
rect 652 31396 692 31436
rect 21772 31312 21812 31352
rect 22636 31312 22676 31352
rect 27916 31312 27956 31352
rect 28780 31312 28820 31352
rect 21388 31228 21428 31268
rect 29164 31228 29204 31268
rect 844 31144 884 31184
rect 23788 31144 23828 31184
rect 26764 31144 26804 31184
rect 4352 30976 4392 31016
rect 4434 30976 4474 31016
rect 4516 30976 4556 31016
rect 4598 30976 4638 31016
rect 4680 30976 4720 31016
rect 19472 30976 19512 31016
rect 19554 30976 19594 31016
rect 19636 30976 19676 31016
rect 19718 30976 19758 31016
rect 19800 30976 19840 31016
rect 34592 30976 34632 31016
rect 34674 30976 34714 31016
rect 34756 30976 34796 31016
rect 34838 30976 34878 31016
rect 34920 30976 34960 31016
rect 49712 30976 49752 31016
rect 49794 30976 49834 31016
rect 49876 30976 49916 31016
rect 49958 30976 49998 31016
rect 50040 30976 50080 31016
rect 64832 30976 64872 31016
rect 64914 30976 64954 31016
rect 64996 30976 65036 31016
rect 65078 30976 65118 31016
rect 65160 30976 65200 31016
rect 79952 30976 79992 31016
rect 80034 30976 80074 31016
rect 80116 30976 80156 31016
rect 80198 30976 80238 31016
rect 80280 30976 80320 31016
rect 95072 30976 95112 31016
rect 95154 30976 95194 31016
rect 95236 30976 95276 31016
rect 95318 30976 95358 31016
rect 95400 30976 95440 31016
rect 27244 30640 27284 30680
rect 27628 30640 27668 30680
rect 32716 30640 32756 30680
rect 33100 30640 33140 30680
rect 33964 30640 34004 30680
rect 652 30556 692 30596
rect 27340 30556 27380 30596
rect 27532 30556 27572 30596
rect 27436 30472 27476 30512
rect 844 30388 884 30428
rect 35116 30388 35156 30428
rect 3112 30220 3152 30260
rect 3194 30220 3234 30260
rect 3276 30220 3316 30260
rect 3358 30220 3398 30260
rect 3440 30220 3480 30260
rect 18232 30220 18272 30260
rect 18314 30220 18354 30260
rect 18396 30220 18436 30260
rect 18478 30220 18518 30260
rect 18560 30220 18600 30260
rect 33352 30220 33392 30260
rect 33434 30220 33474 30260
rect 33516 30220 33556 30260
rect 33598 30220 33638 30260
rect 33680 30220 33720 30260
rect 48472 30220 48512 30260
rect 48554 30220 48594 30260
rect 48636 30220 48676 30260
rect 48718 30220 48758 30260
rect 48800 30220 48840 30260
rect 63592 30220 63632 30260
rect 63674 30220 63714 30260
rect 63756 30220 63796 30260
rect 63838 30220 63878 30260
rect 63920 30220 63960 30260
rect 78712 30220 78752 30260
rect 78794 30220 78834 30260
rect 78876 30220 78916 30260
rect 78958 30220 78998 30260
rect 79040 30220 79080 30260
rect 93832 30220 93872 30260
rect 93914 30220 93954 30260
rect 93996 30220 94036 30260
rect 94078 30220 94118 30260
rect 94160 30220 94200 30260
rect 652 29884 692 29924
rect 36460 29800 36500 29840
rect 844 29632 884 29672
rect 36748 29632 36788 29672
rect 4352 29464 4392 29504
rect 4434 29464 4474 29504
rect 4516 29464 4556 29504
rect 4598 29464 4638 29504
rect 4680 29464 4720 29504
rect 19472 29464 19512 29504
rect 19554 29464 19594 29504
rect 19636 29464 19676 29504
rect 19718 29464 19758 29504
rect 19800 29464 19840 29504
rect 34592 29464 34632 29504
rect 34674 29464 34714 29504
rect 34756 29464 34796 29504
rect 34838 29464 34878 29504
rect 34920 29464 34960 29504
rect 49712 29464 49752 29504
rect 49794 29464 49834 29504
rect 49876 29464 49916 29504
rect 49958 29464 49998 29504
rect 50040 29464 50080 29504
rect 64832 29464 64872 29504
rect 64914 29464 64954 29504
rect 64996 29464 65036 29504
rect 65078 29464 65118 29504
rect 65160 29464 65200 29504
rect 79952 29464 79992 29504
rect 80034 29464 80074 29504
rect 80116 29464 80156 29504
rect 80198 29464 80238 29504
rect 80280 29464 80320 29504
rect 95072 29464 95112 29504
rect 95154 29464 95194 29504
rect 95236 29464 95276 29504
rect 95318 29464 95358 29504
rect 95400 29464 95440 29504
rect 31276 29296 31316 29336
rect 15340 29128 15380 29168
rect 15724 29128 15764 29168
rect 16588 29128 16628 29168
rect 31180 29128 31220 29168
rect 35596 29128 35636 29168
rect 35980 29128 36020 29168
rect 35692 29044 35732 29084
rect 35884 29044 35924 29084
rect 35788 28960 35828 29000
rect 17740 28876 17780 28916
rect 3112 28708 3152 28748
rect 3194 28708 3234 28748
rect 3276 28708 3316 28748
rect 3358 28708 3398 28748
rect 3440 28708 3480 28748
rect 18232 28708 18272 28748
rect 18314 28708 18354 28748
rect 18396 28708 18436 28748
rect 18478 28708 18518 28748
rect 18560 28708 18600 28748
rect 33352 28708 33392 28748
rect 33434 28708 33474 28748
rect 33516 28708 33556 28748
rect 33598 28708 33638 28748
rect 33680 28708 33720 28748
rect 48472 28708 48512 28748
rect 48554 28708 48594 28748
rect 48636 28708 48676 28748
rect 48718 28708 48758 28748
rect 48800 28708 48840 28748
rect 63592 28708 63632 28748
rect 63674 28708 63714 28748
rect 63756 28708 63796 28748
rect 63838 28708 63878 28748
rect 63920 28708 63960 28748
rect 78712 28708 78752 28748
rect 78794 28708 78834 28748
rect 78876 28708 78916 28748
rect 78958 28708 78998 28748
rect 79040 28708 79080 28748
rect 93832 28708 93872 28748
rect 93914 28708 93954 28748
rect 93996 28708 94036 28748
rect 94078 28708 94118 28748
rect 94160 28708 94200 28748
rect 22060 28540 22100 28580
rect 28300 28456 28340 28496
rect 28780 28456 28820 28496
rect 28204 28372 28244 28412
rect 28396 28372 28436 28412
rect 652 28288 692 28328
rect 844 28288 884 28328
rect 22348 28288 22388 28328
rect 22444 28288 22484 28328
rect 23404 28288 23444 28328
rect 28108 28288 28148 28328
rect 28492 28288 28532 28328
rect 29068 28288 29108 28328
rect 29164 28288 29204 28328
rect 29452 28288 29492 28328
rect 29644 28288 29684 28328
rect 29740 28288 29780 28328
rect 23212 28204 23252 28244
rect 23500 28120 23540 28160
rect 29452 28120 29492 28160
rect 22540 28062 22580 28102
rect 29260 28062 29300 28102
rect 4352 27952 4392 27992
rect 4434 27952 4474 27992
rect 4516 27952 4556 27992
rect 4598 27952 4638 27992
rect 4680 27952 4720 27992
rect 19472 27952 19512 27992
rect 19554 27952 19594 27992
rect 19636 27952 19676 27992
rect 19718 27952 19758 27992
rect 19800 27952 19840 27992
rect 34592 27952 34632 27992
rect 34674 27952 34714 27992
rect 34756 27952 34796 27992
rect 34838 27952 34878 27992
rect 34920 27952 34960 27992
rect 49712 27952 49752 27992
rect 49794 27952 49834 27992
rect 49876 27952 49916 27992
rect 49958 27952 49998 27992
rect 50040 27952 50080 27992
rect 64832 27952 64872 27992
rect 64914 27952 64954 27992
rect 64996 27952 65036 27992
rect 65078 27952 65118 27992
rect 65160 27952 65200 27992
rect 79952 27952 79992 27992
rect 80034 27952 80074 27992
rect 80116 27952 80156 27992
rect 80198 27952 80238 27992
rect 80280 27952 80320 27992
rect 95072 27952 95112 27992
rect 95154 27952 95194 27992
rect 95236 27952 95276 27992
rect 95318 27952 95358 27992
rect 95400 27952 95440 27992
rect 20044 27784 20084 27824
rect 23308 27784 23348 27824
rect 26860 27784 26900 27824
rect 26572 27700 26612 27740
rect 27148 27700 27188 27740
rect 652 27616 692 27656
rect 844 27616 884 27656
rect 18124 27616 18164 27656
rect 18508 27616 18548 27656
rect 18700 27616 18740 27656
rect 20140 27616 20180 27656
rect 23404 27616 23444 27656
rect 26380 27616 26420 27656
rect 26668 27616 26708 27656
rect 26956 27616 26996 27656
rect 29548 27616 29588 27656
rect 29644 27600 29684 27640
rect 18220 27532 18260 27572
rect 18412 27532 18452 27572
rect 29452 27532 29492 27572
rect 18316 27448 18356 27488
rect 29260 27448 29300 27488
rect 29356 27406 29396 27446
rect 18796 27364 18836 27404
rect 20332 27364 20372 27404
rect 23596 27364 23636 27404
rect 3112 27196 3152 27236
rect 3194 27196 3234 27236
rect 3276 27196 3316 27236
rect 3358 27196 3398 27236
rect 3440 27196 3480 27236
rect 18232 27196 18272 27236
rect 18314 27196 18354 27236
rect 18396 27196 18436 27236
rect 18478 27196 18518 27236
rect 18560 27196 18600 27236
rect 33352 27196 33392 27236
rect 33434 27196 33474 27236
rect 33516 27196 33556 27236
rect 33598 27196 33638 27236
rect 33680 27196 33720 27236
rect 48472 27196 48512 27236
rect 48554 27196 48594 27236
rect 48636 27196 48676 27236
rect 48718 27196 48758 27236
rect 48800 27196 48840 27236
rect 63592 27196 63632 27236
rect 63674 27196 63714 27236
rect 63756 27196 63796 27236
rect 63838 27196 63878 27236
rect 63920 27196 63960 27236
rect 78712 27196 78752 27236
rect 78794 27196 78834 27236
rect 78876 27196 78916 27236
rect 78958 27196 78998 27236
rect 79040 27196 79080 27236
rect 93832 27196 93872 27236
rect 93914 27196 93954 27236
rect 93996 27196 94036 27236
rect 94078 27196 94118 27236
rect 94160 27196 94200 27236
rect 29452 27028 29492 27068
rect 29932 27028 29972 27068
rect 37324 27028 37364 27068
rect 19948 26944 19988 26984
rect 29644 26944 29684 26984
rect 30124 26944 30164 26984
rect 652 26776 692 26816
rect 844 26776 884 26816
rect 19948 26776 19988 26816
rect 20428 26776 20468 26816
rect 20524 26776 20564 26816
rect 20620 26776 20660 26816
rect 29644 26776 29684 26816
rect 30124 26776 30164 26816
rect 34924 26776 34964 26816
rect 35308 26776 35348 26816
rect 36172 26776 36212 26816
rect 20140 26608 20180 26648
rect 20332 26608 20372 26648
rect 4352 26440 4392 26480
rect 4434 26440 4474 26480
rect 4516 26440 4556 26480
rect 4598 26440 4638 26480
rect 4680 26440 4720 26480
rect 19472 26440 19512 26480
rect 19554 26440 19594 26480
rect 19636 26440 19676 26480
rect 19718 26440 19758 26480
rect 19800 26440 19840 26480
rect 34592 26440 34632 26480
rect 34674 26440 34714 26480
rect 34756 26440 34796 26480
rect 34838 26440 34878 26480
rect 34920 26440 34960 26480
rect 49712 26440 49752 26480
rect 49794 26440 49834 26480
rect 49876 26440 49916 26480
rect 49958 26440 49998 26480
rect 50040 26440 50080 26480
rect 64832 26440 64872 26480
rect 64914 26440 64954 26480
rect 64996 26440 65036 26480
rect 65078 26440 65118 26480
rect 65160 26440 65200 26480
rect 79952 26440 79992 26480
rect 80034 26440 80074 26480
rect 80116 26440 80156 26480
rect 80198 26440 80238 26480
rect 80280 26440 80320 26480
rect 95072 26440 95112 26480
rect 95154 26440 95194 26480
rect 95236 26440 95276 26480
rect 95318 26440 95358 26480
rect 95400 26440 95440 26480
rect 17260 26272 17300 26312
rect 21580 26272 21620 26312
rect 25804 26272 25844 26312
rect 28300 26272 28340 26312
rect 14860 26188 14900 26228
rect 652 26104 692 26144
rect 844 26104 884 26144
rect 15244 26104 15284 26144
rect 16108 26104 16148 26144
rect 21484 26104 21524 26144
rect 21676 26104 21716 26144
rect 21772 26104 21812 26144
rect 26380 26104 26420 26144
rect 27244 26104 27284 26144
rect 28300 26104 28340 26144
rect 28396 26104 28436 26144
rect 34348 26104 34388 26144
rect 35308 26104 35348 26144
rect 39628 26104 39668 26144
rect 25996 26020 26036 26060
rect 28204 26020 28244 26060
rect 28108 25936 28148 25976
rect 39916 25852 39956 25892
rect 3112 25684 3152 25724
rect 3194 25684 3234 25724
rect 3276 25684 3316 25724
rect 3358 25684 3398 25724
rect 3440 25684 3480 25724
rect 18232 25684 18272 25724
rect 18314 25684 18354 25724
rect 18396 25684 18436 25724
rect 18478 25684 18518 25724
rect 18560 25684 18600 25724
rect 33352 25684 33392 25724
rect 33434 25684 33474 25724
rect 33516 25684 33556 25724
rect 33598 25684 33638 25724
rect 33680 25684 33720 25724
rect 48472 25684 48512 25724
rect 48554 25684 48594 25724
rect 48636 25684 48676 25724
rect 48718 25684 48758 25724
rect 48800 25684 48840 25724
rect 63592 25684 63632 25724
rect 63674 25684 63714 25724
rect 63756 25684 63796 25724
rect 63838 25684 63878 25724
rect 63920 25684 63960 25724
rect 78712 25684 78752 25724
rect 78794 25684 78834 25724
rect 78876 25684 78916 25724
rect 78958 25684 78998 25724
rect 79040 25684 79080 25724
rect 93832 25684 93872 25724
rect 93914 25684 93954 25724
rect 93996 25684 94036 25724
rect 94078 25684 94118 25724
rect 94160 25684 94200 25724
rect 28204 25516 28244 25556
rect 652 25264 692 25304
rect 844 25264 884 25304
rect 28396 25264 28436 25304
rect 28492 25096 28532 25136
rect 4352 24928 4392 24968
rect 4434 24928 4474 24968
rect 4516 24928 4556 24968
rect 4598 24928 4638 24968
rect 4680 24928 4720 24968
rect 19472 24928 19512 24968
rect 19554 24928 19594 24968
rect 19636 24928 19676 24968
rect 19718 24928 19758 24968
rect 19800 24928 19840 24968
rect 34592 24928 34632 24968
rect 34674 24928 34714 24968
rect 34756 24928 34796 24968
rect 34838 24928 34878 24968
rect 34920 24928 34960 24968
rect 49712 24928 49752 24968
rect 49794 24928 49834 24968
rect 49876 24928 49916 24968
rect 49958 24928 49998 24968
rect 50040 24928 50080 24968
rect 64832 24928 64872 24968
rect 64914 24928 64954 24968
rect 64996 24928 65036 24968
rect 65078 24928 65118 24968
rect 65160 24928 65200 24968
rect 79952 24928 79992 24968
rect 80034 24928 80074 24968
rect 80116 24928 80156 24968
rect 80198 24928 80238 24968
rect 80280 24928 80320 24968
rect 95072 24928 95112 24968
rect 95154 24928 95194 24968
rect 95236 24928 95276 24968
rect 95318 24928 95358 24968
rect 95400 24928 95440 24968
rect 29644 24760 29684 24800
rect 29836 24676 29876 24716
rect 652 24592 692 24632
rect 844 24592 884 24632
rect 23020 24592 23060 24632
rect 23980 24592 24020 24632
rect 30028 24592 30068 24632
rect 22636 24508 22676 24548
rect 3112 24172 3152 24212
rect 3194 24172 3234 24212
rect 3276 24172 3316 24212
rect 3358 24172 3398 24212
rect 3440 24172 3480 24212
rect 18232 24172 18272 24212
rect 18314 24172 18354 24212
rect 18396 24172 18436 24212
rect 18478 24172 18518 24212
rect 18560 24172 18600 24212
rect 33352 24172 33392 24212
rect 33434 24172 33474 24212
rect 33516 24172 33556 24212
rect 33598 24172 33638 24212
rect 33680 24172 33720 24212
rect 48472 24172 48512 24212
rect 48554 24172 48594 24212
rect 48636 24172 48676 24212
rect 48718 24172 48758 24212
rect 48800 24172 48840 24212
rect 63592 24172 63632 24212
rect 63674 24172 63714 24212
rect 63756 24172 63796 24212
rect 63838 24172 63878 24212
rect 63920 24172 63960 24212
rect 78712 24172 78752 24212
rect 78794 24172 78834 24212
rect 78876 24172 78916 24212
rect 78958 24172 78998 24212
rect 79040 24172 79080 24212
rect 93832 24172 93872 24212
rect 93914 24172 93954 24212
rect 93996 24172 94036 24212
rect 94078 24172 94118 24212
rect 94160 24172 94200 24212
rect 28876 23920 28916 23960
rect 32812 23836 32852 23876
rect 652 23752 692 23792
rect 844 23752 884 23792
rect 28972 23752 29012 23792
rect 33292 23752 33332 23792
rect 33772 23584 33812 23624
rect 4352 23416 4392 23456
rect 4434 23416 4474 23456
rect 4516 23416 4556 23456
rect 4598 23416 4638 23456
rect 4680 23416 4720 23456
rect 19472 23416 19512 23456
rect 19554 23416 19594 23456
rect 19636 23416 19676 23456
rect 19718 23416 19758 23456
rect 19800 23416 19840 23456
rect 34592 23416 34632 23456
rect 34674 23416 34714 23456
rect 34756 23416 34796 23456
rect 34838 23416 34878 23456
rect 34920 23416 34960 23456
rect 49712 23416 49752 23456
rect 49794 23416 49834 23456
rect 49876 23416 49916 23456
rect 49958 23416 49998 23456
rect 50040 23416 50080 23456
rect 64832 23416 64872 23456
rect 64914 23416 64954 23456
rect 64996 23416 65036 23456
rect 65078 23416 65118 23456
rect 65160 23416 65200 23456
rect 79952 23416 79992 23456
rect 80034 23416 80074 23456
rect 80116 23416 80156 23456
rect 80198 23416 80238 23456
rect 80280 23416 80320 23456
rect 95072 23416 95112 23456
rect 95154 23416 95194 23456
rect 95236 23416 95276 23456
rect 95318 23416 95358 23456
rect 95400 23416 95440 23456
rect 19372 23080 19412 23120
rect 19756 23080 19796 23120
rect 20620 23080 20660 23120
rect 28588 23080 28628 23120
rect 28684 23080 28724 23120
rect 28876 23080 28916 23120
rect 34060 23080 34100 23120
rect 34444 23080 34484 23120
rect 35308 23080 35348 23120
rect 21772 22828 21812 22868
rect 28876 22828 28916 22868
rect 36460 22828 36500 22868
rect 3112 22660 3152 22700
rect 3194 22660 3234 22700
rect 3276 22660 3316 22700
rect 3358 22660 3398 22700
rect 3440 22660 3480 22700
rect 18232 22660 18272 22700
rect 18314 22660 18354 22700
rect 18396 22660 18436 22700
rect 18478 22660 18518 22700
rect 18560 22660 18600 22700
rect 33352 22660 33392 22700
rect 33434 22660 33474 22700
rect 33516 22660 33556 22700
rect 33598 22660 33638 22700
rect 33680 22660 33720 22700
rect 48472 22660 48512 22700
rect 48554 22660 48594 22700
rect 48636 22660 48676 22700
rect 48718 22660 48758 22700
rect 48800 22660 48840 22700
rect 63592 22660 63632 22700
rect 63674 22660 63714 22700
rect 63756 22660 63796 22700
rect 63838 22660 63878 22700
rect 63920 22660 63960 22700
rect 78712 22660 78752 22700
rect 78794 22660 78834 22700
rect 78876 22660 78916 22700
rect 78958 22660 78998 22700
rect 79040 22660 79080 22700
rect 93832 22660 93872 22700
rect 93914 22660 93954 22700
rect 93996 22660 94036 22700
rect 94078 22660 94118 22700
rect 94160 22660 94200 22700
rect 652 22408 692 22448
rect 29164 22408 29204 22448
rect 26572 22324 26612 22364
rect 35308 22324 35348 22364
rect 41548 22324 41588 22364
rect 15340 22240 15380 22280
rect 16204 22240 16244 22280
rect 24556 22240 24596 22280
rect 25420 22240 25460 22280
rect 28684 22240 28724 22280
rect 28780 22240 28820 22280
rect 28876 22240 28916 22280
rect 29260 22240 29300 22280
rect 32428 22240 32468 22280
rect 32524 22240 32564 22280
rect 32620 22240 32660 22280
rect 34060 22240 34100 22280
rect 34156 22240 34196 22280
rect 34924 22240 34964 22280
rect 35020 22240 35060 22280
rect 35212 22240 35252 22280
rect 35404 22240 35444 22280
rect 35596 22240 35636 22280
rect 35788 22240 35828 22280
rect 39532 22240 39572 22280
rect 40396 22240 40436 22280
rect 14956 22156 14996 22196
rect 24172 22156 24212 22196
rect 34252 22156 34292 22196
rect 34820 22156 34860 22196
rect 35692 22156 35732 22196
rect 39148 22156 39188 22196
rect 17356 22072 17396 22112
rect 28972 22072 29012 22112
rect 34348 22072 34388 22112
rect 34444 22072 34484 22112
rect 34636 22072 34676 22112
rect 34732 22072 34772 22112
rect 4352 21904 4392 21944
rect 4434 21904 4474 21944
rect 4516 21904 4556 21944
rect 4598 21904 4638 21944
rect 4680 21904 4720 21944
rect 19472 21904 19512 21944
rect 19554 21904 19594 21944
rect 19636 21904 19676 21944
rect 19718 21904 19758 21944
rect 19800 21904 19840 21944
rect 34592 21904 34632 21944
rect 34674 21904 34714 21944
rect 34756 21904 34796 21944
rect 34838 21904 34878 21944
rect 34920 21904 34960 21944
rect 49712 21904 49752 21944
rect 49794 21904 49834 21944
rect 49876 21904 49916 21944
rect 49958 21904 49998 21944
rect 50040 21904 50080 21944
rect 64832 21904 64872 21944
rect 64914 21904 64954 21944
rect 64996 21904 65036 21944
rect 65078 21904 65118 21944
rect 65160 21904 65200 21944
rect 79952 21904 79992 21944
rect 80034 21904 80074 21944
rect 80116 21904 80156 21944
rect 80198 21904 80238 21944
rect 80280 21904 80320 21944
rect 95072 21904 95112 21944
rect 95154 21904 95194 21944
rect 95236 21904 95276 21944
rect 95318 21904 95358 21944
rect 95400 21904 95440 21944
rect 28396 21568 28436 21608
rect 29356 21568 29396 21608
rect 3112 21148 3152 21188
rect 3194 21148 3234 21188
rect 3276 21148 3316 21188
rect 3358 21148 3398 21188
rect 3440 21148 3480 21188
rect 18232 21148 18272 21188
rect 18314 21148 18354 21188
rect 18396 21148 18436 21188
rect 18478 21148 18518 21188
rect 18560 21148 18600 21188
rect 33352 21148 33392 21188
rect 33434 21148 33474 21188
rect 33516 21148 33556 21188
rect 33598 21148 33638 21188
rect 33680 21148 33720 21188
rect 48472 21148 48512 21188
rect 48554 21148 48594 21188
rect 48636 21148 48676 21188
rect 48718 21148 48758 21188
rect 48800 21148 48840 21188
rect 63592 21148 63632 21188
rect 63674 21148 63714 21188
rect 63756 21148 63796 21188
rect 63838 21148 63878 21188
rect 63920 21148 63960 21188
rect 78712 21148 78752 21188
rect 78794 21148 78834 21188
rect 78876 21148 78916 21188
rect 78958 21148 78998 21188
rect 79040 21148 79080 21188
rect 93832 21148 93872 21188
rect 93914 21148 93954 21188
rect 93996 21148 94036 21188
rect 94078 21148 94118 21188
rect 94160 21148 94200 21188
rect 19180 20980 19220 21020
rect 652 20896 692 20936
rect 30604 20896 30644 20936
rect 30796 20812 30836 20852
rect 31372 20812 31412 20852
rect 19372 20728 19412 20768
rect 19468 20728 19508 20768
rect 19564 20728 19604 20768
rect 22636 20728 22676 20768
rect 22732 20728 22772 20768
rect 22828 20728 22868 20768
rect 23116 20728 23156 20768
rect 23212 20728 23252 20768
rect 23308 20728 23348 20768
rect 23404 20728 23444 20768
rect 29164 20728 29204 20768
rect 30316 20728 30356 20768
rect 30508 20728 30548 20768
rect 30604 20728 30644 20768
rect 31180 20728 31220 20768
rect 22924 20644 22964 20684
rect 29452 20560 29492 20600
rect 29644 20560 29684 20600
rect 30892 20560 30932 20600
rect 4352 20392 4392 20432
rect 4434 20392 4474 20432
rect 4516 20392 4556 20432
rect 4598 20392 4638 20432
rect 4680 20392 4720 20432
rect 19472 20392 19512 20432
rect 19554 20392 19594 20432
rect 19636 20392 19676 20432
rect 19718 20392 19758 20432
rect 19800 20392 19840 20432
rect 34592 20392 34632 20432
rect 34674 20392 34714 20432
rect 34756 20392 34796 20432
rect 34838 20392 34878 20432
rect 34920 20392 34960 20432
rect 49712 20392 49752 20432
rect 49794 20392 49834 20432
rect 49876 20392 49916 20432
rect 49958 20392 49998 20432
rect 50040 20392 50080 20432
rect 64832 20392 64872 20432
rect 64914 20392 64954 20432
rect 64996 20392 65036 20432
rect 65078 20392 65118 20432
rect 65160 20392 65200 20432
rect 79952 20392 79992 20432
rect 80034 20392 80074 20432
rect 80116 20392 80156 20432
rect 80198 20392 80238 20432
rect 80280 20392 80320 20432
rect 95072 20392 95112 20432
rect 95154 20392 95194 20432
rect 95236 20392 95276 20432
rect 95318 20392 95358 20432
rect 95400 20392 95440 20432
rect 22060 20224 22100 20264
rect 15436 20140 15476 20180
rect 34924 20140 34964 20180
rect 15628 20056 15668 20096
rect 15916 20056 15956 20096
rect 21100 20056 21140 20096
rect 21196 20056 21236 20096
rect 21388 20056 21428 20096
rect 21772 20056 21812 20096
rect 21868 20056 21908 20096
rect 23212 20056 23252 20096
rect 24172 20056 24212 20096
rect 34828 20056 34868 20096
rect 35020 20056 35060 20096
rect 39916 20056 39956 20096
rect 22828 19972 22868 20012
rect 652 19888 692 19928
rect 21388 19888 21428 19928
rect 23692 19804 23732 19844
rect 39244 19804 39284 19844
rect 3112 19636 3152 19676
rect 3194 19636 3234 19676
rect 3276 19636 3316 19676
rect 3358 19636 3398 19676
rect 3440 19636 3480 19676
rect 18232 19636 18272 19676
rect 18314 19636 18354 19676
rect 18396 19636 18436 19676
rect 18478 19636 18518 19676
rect 18560 19636 18600 19676
rect 33352 19636 33392 19676
rect 33434 19636 33474 19676
rect 33516 19636 33556 19676
rect 33598 19636 33638 19676
rect 33680 19636 33720 19676
rect 48472 19636 48512 19676
rect 48554 19636 48594 19676
rect 48636 19636 48676 19676
rect 48718 19636 48758 19676
rect 48800 19636 48840 19676
rect 63592 19636 63632 19676
rect 63674 19636 63714 19676
rect 63756 19636 63796 19676
rect 63838 19636 63878 19676
rect 63920 19636 63960 19676
rect 78712 19636 78752 19676
rect 78794 19636 78834 19676
rect 78876 19636 78916 19676
rect 78958 19636 78998 19676
rect 79040 19636 79080 19676
rect 93832 19636 93872 19676
rect 93914 19636 93954 19676
rect 93996 19636 94036 19676
rect 94078 19636 94118 19676
rect 94160 19636 94200 19676
rect 41164 19468 41204 19508
rect 652 19384 692 19424
rect 33868 19384 33908 19424
rect 37516 19384 37556 19424
rect 19180 19300 19220 19340
rect 19084 19216 19124 19256
rect 19468 19216 19508 19256
rect 19660 19216 19700 19256
rect 33196 19216 33236 19256
rect 36844 19216 36884 19256
rect 37132 19216 37172 19256
rect 37228 19216 37268 19256
rect 38764 19216 38804 19256
rect 39148 19216 39188 19256
rect 40012 19216 40052 19256
rect 19468 19048 19508 19088
rect 4352 18880 4392 18920
rect 4434 18880 4474 18920
rect 4516 18880 4556 18920
rect 4598 18880 4638 18920
rect 4680 18880 4720 18920
rect 19472 18880 19512 18920
rect 19554 18880 19594 18920
rect 19636 18880 19676 18920
rect 19718 18880 19758 18920
rect 19800 18880 19840 18920
rect 34592 18880 34632 18920
rect 34674 18880 34714 18920
rect 34756 18880 34796 18920
rect 34838 18880 34878 18920
rect 34920 18880 34960 18920
rect 49712 18880 49752 18920
rect 49794 18880 49834 18920
rect 49876 18880 49916 18920
rect 49958 18880 49998 18920
rect 50040 18880 50080 18920
rect 64832 18880 64872 18920
rect 64914 18880 64954 18920
rect 64996 18880 65036 18920
rect 65078 18880 65118 18920
rect 65160 18880 65200 18920
rect 79952 18880 79992 18920
rect 80034 18880 80074 18920
rect 80116 18880 80156 18920
rect 80198 18880 80238 18920
rect 80280 18880 80320 18920
rect 95072 18880 95112 18920
rect 95154 18880 95194 18920
rect 95236 18880 95276 18920
rect 95318 18880 95358 18920
rect 95400 18880 95440 18920
rect 17548 18628 17588 18668
rect 27340 18628 27380 18668
rect 17740 18544 17780 18584
rect 18028 18544 18068 18584
rect 22444 18544 22484 18584
rect 26092 18544 26132 18584
rect 26476 18544 26516 18584
rect 27436 18544 27476 18584
rect 28396 18544 28436 18584
rect 29068 18544 29108 18584
rect 22252 18460 22292 18500
rect 26188 18460 26228 18500
rect 26380 18460 26420 18500
rect 652 18376 692 18416
rect 26284 18376 26324 18416
rect 22444 18292 22484 18332
rect 3112 18124 3152 18164
rect 3194 18124 3234 18164
rect 3276 18124 3316 18164
rect 3358 18124 3398 18164
rect 3440 18124 3480 18164
rect 18232 18124 18272 18164
rect 18314 18124 18354 18164
rect 18396 18124 18436 18164
rect 18478 18124 18518 18164
rect 18560 18124 18600 18164
rect 33352 18124 33392 18164
rect 33434 18124 33474 18164
rect 33516 18124 33556 18164
rect 33598 18124 33638 18164
rect 33680 18124 33720 18164
rect 48472 18124 48512 18164
rect 48554 18124 48594 18164
rect 48636 18124 48676 18164
rect 48718 18124 48758 18164
rect 48800 18124 48840 18164
rect 63592 18124 63632 18164
rect 63674 18124 63714 18164
rect 63756 18124 63796 18164
rect 63838 18124 63878 18164
rect 63920 18124 63960 18164
rect 78712 18124 78752 18164
rect 78794 18124 78834 18164
rect 78876 18124 78916 18164
rect 78958 18124 78998 18164
rect 79040 18124 79080 18164
rect 93832 18124 93872 18164
rect 93914 18124 93954 18164
rect 93996 18124 94036 18164
rect 94078 18124 94118 18164
rect 94160 18124 94200 18164
rect 21388 17956 21428 17996
rect 21868 17956 21908 17996
rect 652 17872 692 17912
rect 22828 17872 22868 17912
rect 29164 17788 29204 17828
rect 16108 17704 16148 17744
rect 16204 17704 16244 17744
rect 21292 17704 21332 17744
rect 21772 17704 21812 17744
rect 22156 17704 22196 17744
rect 22348 17704 22388 17744
rect 22540 17704 22580 17744
rect 22732 17704 22772 17744
rect 22828 17704 22868 17744
rect 26764 17704 26804 17744
rect 27148 17704 27188 17744
rect 28012 17704 28052 17744
rect 33676 17704 33716 17744
rect 33868 17704 33908 17744
rect 37900 17704 37940 17744
rect 38764 17704 38804 17744
rect 22252 17620 22292 17660
rect 33772 17620 33812 17660
rect 15820 17536 15860 17576
rect 4352 17368 4392 17408
rect 4434 17368 4474 17408
rect 4516 17368 4556 17408
rect 4598 17368 4638 17408
rect 4680 17368 4720 17408
rect 19472 17368 19512 17408
rect 19554 17368 19594 17408
rect 19636 17368 19676 17408
rect 19718 17368 19758 17408
rect 19800 17368 19840 17408
rect 34592 17368 34632 17408
rect 34674 17368 34714 17408
rect 34756 17368 34796 17408
rect 34838 17368 34878 17408
rect 34920 17368 34960 17408
rect 49712 17368 49752 17408
rect 49794 17368 49834 17408
rect 49876 17368 49916 17408
rect 49958 17368 49998 17408
rect 50040 17368 50080 17408
rect 64832 17368 64872 17408
rect 64914 17368 64954 17408
rect 64996 17368 65036 17408
rect 65078 17368 65118 17408
rect 65160 17368 65200 17408
rect 79952 17368 79992 17408
rect 80034 17368 80074 17408
rect 80116 17368 80156 17408
rect 80198 17368 80238 17408
rect 80280 17368 80320 17408
rect 95072 17368 95112 17408
rect 95154 17368 95194 17408
rect 95236 17368 95276 17408
rect 95318 17368 95358 17408
rect 95400 17368 95440 17408
rect 31372 17116 31412 17156
rect 15820 17032 15860 17072
rect 16012 17032 16052 17072
rect 22060 17032 22100 17072
rect 22252 17032 22292 17072
rect 22348 17032 22388 17072
rect 31756 17032 31796 17072
rect 32620 17032 32660 17072
rect 34252 17032 34292 17072
rect 15916 16948 15956 16988
rect 33772 16948 33812 16988
rect 34060 16948 34100 16988
rect 652 16864 692 16904
rect 22348 16864 22388 16904
rect 34252 16780 34292 16820
rect 3112 16612 3152 16652
rect 3194 16612 3234 16652
rect 3276 16612 3316 16652
rect 3358 16612 3398 16652
rect 3440 16612 3480 16652
rect 18232 16612 18272 16652
rect 18314 16612 18354 16652
rect 18396 16612 18436 16652
rect 18478 16612 18518 16652
rect 18560 16612 18600 16652
rect 33352 16612 33392 16652
rect 33434 16612 33474 16652
rect 33516 16612 33556 16652
rect 33598 16612 33638 16652
rect 33680 16612 33720 16652
rect 48472 16612 48512 16652
rect 48554 16612 48594 16652
rect 48636 16612 48676 16652
rect 48718 16612 48758 16652
rect 48800 16612 48840 16652
rect 63592 16612 63632 16652
rect 63674 16612 63714 16652
rect 63756 16612 63796 16652
rect 63838 16612 63878 16652
rect 63920 16612 63960 16652
rect 78712 16612 78752 16652
rect 78794 16612 78834 16652
rect 78876 16612 78916 16652
rect 78958 16612 78998 16652
rect 79040 16612 79080 16652
rect 93832 16612 93872 16652
rect 93914 16612 93954 16652
rect 93996 16612 94036 16652
rect 94078 16612 94118 16652
rect 94160 16612 94200 16652
rect 652 16360 692 16400
rect 33964 16360 34004 16400
rect 33868 16276 33908 16316
rect 34060 16276 34100 16316
rect 33772 16192 33812 16232
rect 34156 16192 34196 16232
rect 37228 16192 37268 16232
rect 37324 16192 37364 16232
rect 38572 16192 38612 16232
rect 39244 16192 39284 16232
rect 37036 16024 37076 16064
rect 4352 15856 4392 15896
rect 4434 15856 4474 15896
rect 4516 15856 4556 15896
rect 4598 15856 4638 15896
rect 4680 15856 4720 15896
rect 19472 15856 19512 15896
rect 19554 15856 19594 15896
rect 19636 15856 19676 15896
rect 19718 15856 19758 15896
rect 19800 15856 19840 15896
rect 34592 15856 34632 15896
rect 34674 15856 34714 15896
rect 34756 15856 34796 15896
rect 34838 15856 34878 15896
rect 34920 15856 34960 15896
rect 49712 15856 49752 15896
rect 49794 15856 49834 15896
rect 49876 15856 49916 15896
rect 49958 15856 49998 15896
rect 50040 15856 50080 15896
rect 64832 15856 64872 15896
rect 64914 15856 64954 15896
rect 64996 15856 65036 15896
rect 65078 15856 65118 15896
rect 65160 15856 65200 15896
rect 79952 15856 79992 15896
rect 80034 15856 80074 15896
rect 80116 15856 80156 15896
rect 80198 15856 80238 15896
rect 80280 15856 80320 15896
rect 95072 15856 95112 15896
rect 95154 15856 95194 15896
rect 95236 15856 95276 15896
rect 95318 15856 95358 15896
rect 95400 15856 95440 15896
rect 652 15688 692 15728
rect 17836 15688 17876 15728
rect 18220 15688 18260 15728
rect 40012 15688 40052 15728
rect 15436 15604 15476 15644
rect 37612 15604 37652 15644
rect 15820 15520 15860 15560
rect 16684 15520 16724 15560
rect 18316 15520 18356 15560
rect 27916 15520 27956 15560
rect 28300 15520 28340 15560
rect 37996 15520 38036 15560
rect 38860 15520 38900 15560
rect 18892 15436 18932 15476
rect 28012 15436 28052 15476
rect 28204 15436 28244 15476
rect 18508 15352 18548 15392
rect 28108 15352 28148 15392
rect 18700 15268 18740 15308
rect 3112 15100 3152 15140
rect 3194 15100 3234 15140
rect 3276 15100 3316 15140
rect 3358 15100 3398 15140
rect 3440 15100 3480 15140
rect 18232 15100 18272 15140
rect 18314 15100 18354 15140
rect 18396 15100 18436 15140
rect 18478 15100 18518 15140
rect 18560 15100 18600 15140
rect 33352 15100 33392 15140
rect 33434 15100 33474 15140
rect 33516 15100 33556 15140
rect 33598 15100 33638 15140
rect 33680 15100 33720 15140
rect 48472 15100 48512 15140
rect 48554 15100 48594 15140
rect 48636 15100 48676 15140
rect 48718 15100 48758 15140
rect 48800 15100 48840 15140
rect 63592 15100 63632 15140
rect 63674 15100 63714 15140
rect 63756 15100 63796 15140
rect 63838 15100 63878 15140
rect 63920 15100 63960 15140
rect 78712 15100 78752 15140
rect 78794 15100 78834 15140
rect 78876 15100 78916 15140
rect 78958 15100 78998 15140
rect 79040 15100 79080 15140
rect 93832 15100 93872 15140
rect 93914 15100 93954 15140
rect 93996 15100 94036 15140
rect 94078 15100 94118 15140
rect 94160 15100 94200 15140
rect 25036 14932 25076 14972
rect 22636 14680 22676 14720
rect 23020 14680 23060 14720
rect 23884 14680 23924 14720
rect 652 14512 692 14552
rect 4352 14344 4392 14384
rect 4434 14344 4474 14384
rect 4516 14344 4556 14384
rect 4598 14344 4638 14384
rect 4680 14344 4720 14384
rect 19472 14344 19512 14384
rect 19554 14344 19594 14384
rect 19636 14344 19676 14384
rect 19718 14344 19758 14384
rect 19800 14344 19840 14384
rect 34592 14344 34632 14384
rect 34674 14344 34714 14384
rect 34756 14344 34796 14384
rect 34838 14344 34878 14384
rect 34920 14344 34960 14384
rect 49712 14344 49752 14384
rect 49794 14344 49834 14384
rect 49876 14344 49916 14384
rect 49958 14344 49998 14384
rect 50040 14344 50080 14384
rect 64832 14344 64872 14384
rect 64914 14344 64954 14384
rect 64996 14344 65036 14384
rect 65078 14344 65118 14384
rect 65160 14344 65200 14384
rect 79952 14344 79992 14384
rect 80034 14344 80074 14384
rect 80116 14344 80156 14384
rect 80198 14344 80238 14384
rect 80280 14344 80320 14384
rect 95072 14344 95112 14384
rect 95154 14344 95194 14384
rect 95236 14344 95276 14384
rect 95318 14344 95358 14384
rect 95400 14344 95440 14384
rect 3112 13588 3152 13628
rect 3194 13588 3234 13628
rect 3276 13588 3316 13628
rect 3358 13588 3398 13628
rect 3440 13588 3480 13628
rect 18232 13588 18272 13628
rect 18314 13588 18354 13628
rect 18396 13588 18436 13628
rect 18478 13588 18518 13628
rect 18560 13588 18600 13628
rect 33352 13588 33392 13628
rect 33434 13588 33474 13628
rect 33516 13588 33556 13628
rect 33598 13588 33638 13628
rect 33680 13588 33720 13628
rect 48472 13588 48512 13628
rect 48554 13588 48594 13628
rect 48636 13588 48676 13628
rect 48718 13588 48758 13628
rect 48800 13588 48840 13628
rect 63592 13588 63632 13628
rect 63674 13588 63714 13628
rect 63756 13588 63796 13628
rect 63838 13588 63878 13628
rect 63920 13588 63960 13628
rect 78712 13588 78752 13628
rect 78794 13588 78834 13628
rect 78876 13588 78916 13628
rect 78958 13588 78998 13628
rect 79040 13588 79080 13628
rect 93832 13588 93872 13628
rect 93914 13588 93954 13628
rect 93996 13588 94036 13628
rect 94078 13588 94118 13628
rect 94160 13588 94200 13628
rect 33196 13168 33236 13208
rect 652 13000 692 13040
rect 33004 13000 33044 13040
rect 33292 13000 33332 13040
rect 4352 12832 4392 12872
rect 4434 12832 4474 12872
rect 4516 12832 4556 12872
rect 4598 12832 4638 12872
rect 4680 12832 4720 12872
rect 19472 12832 19512 12872
rect 19554 12832 19594 12872
rect 19636 12832 19676 12872
rect 19718 12832 19758 12872
rect 19800 12832 19840 12872
rect 34592 12832 34632 12872
rect 34674 12832 34714 12872
rect 34756 12832 34796 12872
rect 34838 12832 34878 12872
rect 34920 12832 34960 12872
rect 49712 12832 49752 12872
rect 49794 12832 49834 12872
rect 49876 12832 49916 12872
rect 49958 12832 49998 12872
rect 50040 12832 50080 12872
rect 64832 12832 64872 12872
rect 64914 12832 64954 12872
rect 64996 12832 65036 12872
rect 65078 12832 65118 12872
rect 65160 12832 65200 12872
rect 79952 12832 79992 12872
rect 80034 12832 80074 12872
rect 80116 12832 80156 12872
rect 80198 12832 80238 12872
rect 80280 12832 80320 12872
rect 95072 12832 95112 12872
rect 95154 12832 95194 12872
rect 95236 12832 95276 12872
rect 95318 12832 95358 12872
rect 95400 12832 95440 12872
rect 652 12664 692 12704
rect 17740 12580 17780 12620
rect 26476 12580 26516 12620
rect 26860 12580 26900 12620
rect 18124 12496 18164 12536
rect 18988 12496 19028 12536
rect 26380 12496 26420 12536
rect 26572 12496 26612 12536
rect 26764 12496 26804 12536
rect 26956 12496 26996 12536
rect 27244 12496 27284 12536
rect 27820 12496 27860 12536
rect 30892 12496 30932 12536
rect 31276 12496 31316 12536
rect 32140 12496 32180 12536
rect 33292 12496 33332 12536
rect 27436 12412 27476 12452
rect 28012 12412 28052 12452
rect 30700 12328 30740 12368
rect 20140 12244 20180 12284
rect 27244 12244 27284 12284
rect 27820 12244 27860 12284
rect 3112 12076 3152 12116
rect 3194 12076 3234 12116
rect 3276 12076 3316 12116
rect 3358 12076 3398 12116
rect 3440 12076 3480 12116
rect 18232 12076 18272 12116
rect 18314 12076 18354 12116
rect 18396 12076 18436 12116
rect 18478 12076 18518 12116
rect 18560 12076 18600 12116
rect 33352 12076 33392 12116
rect 33434 12076 33474 12116
rect 33516 12076 33556 12116
rect 33598 12076 33638 12116
rect 33680 12076 33720 12116
rect 48472 12076 48512 12116
rect 48554 12076 48594 12116
rect 48636 12076 48676 12116
rect 48718 12076 48758 12116
rect 48800 12076 48840 12116
rect 63592 12076 63632 12116
rect 63674 12076 63714 12116
rect 63756 12076 63796 12116
rect 63838 12076 63878 12116
rect 63920 12076 63960 12116
rect 78712 12076 78752 12116
rect 78794 12076 78834 12116
rect 78876 12076 78916 12116
rect 78958 12076 78998 12116
rect 79040 12076 79080 12116
rect 93832 12076 93872 12116
rect 93914 12076 93954 12116
rect 93996 12076 94036 12116
rect 94078 12076 94118 12116
rect 94160 12076 94200 12116
rect 24940 11908 24980 11948
rect 844 11740 884 11780
rect 22540 11656 22580 11696
rect 22924 11656 22964 11696
rect 23788 11656 23828 11696
rect 652 11488 692 11528
rect 4352 11320 4392 11360
rect 4434 11320 4474 11360
rect 4516 11320 4556 11360
rect 4598 11320 4638 11360
rect 4680 11320 4720 11360
rect 19472 11320 19512 11360
rect 19554 11320 19594 11360
rect 19636 11320 19676 11360
rect 19718 11320 19758 11360
rect 19800 11320 19840 11360
rect 34592 11320 34632 11360
rect 34674 11320 34714 11360
rect 34756 11320 34796 11360
rect 34838 11320 34878 11360
rect 34920 11320 34960 11360
rect 49712 11320 49752 11360
rect 49794 11320 49834 11360
rect 49876 11320 49916 11360
rect 49958 11320 49998 11360
rect 50040 11320 50080 11360
rect 64832 11320 64872 11360
rect 64914 11320 64954 11360
rect 64996 11320 65036 11360
rect 65078 11320 65118 11360
rect 65160 11320 65200 11360
rect 79952 11320 79992 11360
rect 80034 11320 80074 11360
rect 80116 11320 80156 11360
rect 80198 11320 80238 11360
rect 80280 11320 80320 11360
rect 95072 11320 95112 11360
rect 95154 11320 95194 11360
rect 95236 11320 95276 11360
rect 95318 11320 95358 11360
rect 95400 11320 95440 11360
rect 844 10900 884 10940
rect 652 10732 692 10772
rect 3112 10564 3152 10604
rect 3194 10564 3234 10604
rect 3276 10564 3316 10604
rect 3358 10564 3398 10604
rect 3440 10564 3480 10604
rect 18232 10564 18272 10604
rect 18314 10564 18354 10604
rect 18396 10564 18436 10604
rect 18478 10564 18518 10604
rect 18560 10564 18600 10604
rect 33352 10564 33392 10604
rect 33434 10564 33474 10604
rect 33516 10564 33556 10604
rect 33598 10564 33638 10604
rect 33680 10564 33720 10604
rect 48472 10564 48512 10604
rect 48554 10564 48594 10604
rect 48636 10564 48676 10604
rect 48718 10564 48758 10604
rect 48800 10564 48840 10604
rect 63592 10564 63632 10604
rect 63674 10564 63714 10604
rect 63756 10564 63796 10604
rect 63838 10564 63878 10604
rect 63920 10564 63960 10604
rect 78712 10564 78752 10604
rect 78794 10564 78834 10604
rect 78876 10564 78916 10604
rect 78958 10564 78998 10604
rect 79040 10564 79080 10604
rect 93832 10564 93872 10604
rect 93914 10564 93954 10604
rect 93996 10564 94036 10604
rect 94078 10564 94118 10604
rect 94160 10564 94200 10604
rect 844 10228 884 10268
rect 652 9976 692 10016
rect 4352 9808 4392 9848
rect 4434 9808 4474 9848
rect 4516 9808 4556 9848
rect 4598 9808 4638 9848
rect 4680 9808 4720 9848
rect 19472 9808 19512 9848
rect 19554 9808 19594 9848
rect 19636 9808 19676 9848
rect 19718 9808 19758 9848
rect 19800 9808 19840 9848
rect 34592 9808 34632 9848
rect 34674 9808 34714 9848
rect 34756 9808 34796 9848
rect 34838 9808 34878 9848
rect 34920 9808 34960 9848
rect 49712 9808 49752 9848
rect 49794 9808 49834 9848
rect 49876 9808 49916 9848
rect 49958 9808 49998 9848
rect 50040 9808 50080 9848
rect 64832 9808 64872 9848
rect 64914 9808 64954 9848
rect 64996 9808 65036 9848
rect 65078 9808 65118 9848
rect 65160 9808 65200 9848
rect 79952 9808 79992 9848
rect 80034 9808 80074 9848
rect 80116 9808 80156 9848
rect 80198 9808 80238 9848
rect 80280 9808 80320 9848
rect 95072 9808 95112 9848
rect 95154 9808 95194 9848
rect 95236 9808 95276 9848
rect 95318 9808 95358 9848
rect 95400 9808 95440 9848
rect 844 9388 884 9428
rect 652 9220 692 9260
rect 3112 9052 3152 9092
rect 3194 9052 3234 9092
rect 3276 9052 3316 9092
rect 3358 9052 3398 9092
rect 3440 9052 3480 9092
rect 18232 9052 18272 9092
rect 18314 9052 18354 9092
rect 18396 9052 18436 9092
rect 18478 9052 18518 9092
rect 18560 9052 18600 9092
rect 33352 9052 33392 9092
rect 33434 9052 33474 9092
rect 33516 9052 33556 9092
rect 33598 9052 33638 9092
rect 33680 9052 33720 9092
rect 48472 9052 48512 9092
rect 48554 9052 48594 9092
rect 48636 9052 48676 9092
rect 48718 9052 48758 9092
rect 48800 9052 48840 9092
rect 63592 9052 63632 9092
rect 63674 9052 63714 9092
rect 63756 9052 63796 9092
rect 63838 9052 63878 9092
rect 63920 9052 63960 9092
rect 78712 9052 78752 9092
rect 78794 9052 78834 9092
rect 78876 9052 78916 9092
rect 78958 9052 78998 9092
rect 79040 9052 79080 9092
rect 93832 9052 93872 9092
rect 93914 9052 93954 9092
rect 93996 9052 94036 9092
rect 94078 9052 94118 9092
rect 94160 9052 94200 9092
rect 844 8716 884 8756
rect 652 8464 692 8504
rect 4352 8296 4392 8336
rect 4434 8296 4474 8336
rect 4516 8296 4556 8336
rect 4598 8296 4638 8336
rect 4680 8296 4720 8336
rect 19472 8296 19512 8336
rect 19554 8296 19594 8336
rect 19636 8296 19676 8336
rect 19718 8296 19758 8336
rect 19800 8296 19840 8336
rect 34592 8296 34632 8336
rect 34674 8296 34714 8336
rect 34756 8296 34796 8336
rect 34838 8296 34878 8336
rect 34920 8296 34960 8336
rect 49712 8296 49752 8336
rect 49794 8296 49834 8336
rect 49876 8296 49916 8336
rect 49958 8296 49998 8336
rect 50040 8296 50080 8336
rect 64832 8296 64872 8336
rect 64914 8296 64954 8336
rect 64996 8296 65036 8336
rect 65078 8296 65118 8336
rect 65160 8296 65200 8336
rect 79952 8296 79992 8336
rect 80034 8296 80074 8336
rect 80116 8296 80156 8336
rect 80198 8296 80238 8336
rect 80280 8296 80320 8336
rect 95072 8296 95112 8336
rect 95154 8296 95194 8336
rect 95236 8296 95276 8336
rect 95318 8296 95358 8336
rect 95400 8296 95440 8336
rect 844 7876 884 7916
rect 652 7708 692 7748
rect 3112 7540 3152 7580
rect 3194 7540 3234 7580
rect 3276 7540 3316 7580
rect 3358 7540 3398 7580
rect 3440 7540 3480 7580
rect 18232 7540 18272 7580
rect 18314 7540 18354 7580
rect 18396 7540 18436 7580
rect 18478 7540 18518 7580
rect 18560 7540 18600 7580
rect 33352 7540 33392 7580
rect 33434 7540 33474 7580
rect 33516 7540 33556 7580
rect 33598 7540 33638 7580
rect 33680 7540 33720 7580
rect 48472 7540 48512 7580
rect 48554 7540 48594 7580
rect 48636 7540 48676 7580
rect 48718 7540 48758 7580
rect 48800 7540 48840 7580
rect 63592 7540 63632 7580
rect 63674 7540 63714 7580
rect 63756 7540 63796 7580
rect 63838 7540 63878 7580
rect 63920 7540 63960 7580
rect 78712 7540 78752 7580
rect 78794 7540 78834 7580
rect 78876 7540 78916 7580
rect 78958 7540 78998 7580
rect 79040 7540 79080 7580
rect 93832 7540 93872 7580
rect 93914 7540 93954 7580
rect 93996 7540 94036 7580
rect 94078 7540 94118 7580
rect 94160 7540 94200 7580
rect 844 7204 884 7244
rect 652 6952 692 6992
rect 4352 6784 4392 6824
rect 4434 6784 4474 6824
rect 4516 6784 4556 6824
rect 4598 6784 4638 6824
rect 4680 6784 4720 6824
rect 19472 6784 19512 6824
rect 19554 6784 19594 6824
rect 19636 6784 19676 6824
rect 19718 6784 19758 6824
rect 19800 6784 19840 6824
rect 34592 6784 34632 6824
rect 34674 6784 34714 6824
rect 34756 6784 34796 6824
rect 34838 6784 34878 6824
rect 34920 6784 34960 6824
rect 49712 6784 49752 6824
rect 49794 6784 49834 6824
rect 49876 6784 49916 6824
rect 49958 6784 49998 6824
rect 50040 6784 50080 6824
rect 64832 6784 64872 6824
rect 64914 6784 64954 6824
rect 64996 6784 65036 6824
rect 65078 6784 65118 6824
rect 65160 6784 65200 6824
rect 79952 6784 79992 6824
rect 80034 6784 80074 6824
rect 80116 6784 80156 6824
rect 80198 6784 80238 6824
rect 80280 6784 80320 6824
rect 95072 6784 95112 6824
rect 95154 6784 95194 6824
rect 95236 6784 95276 6824
rect 95318 6784 95358 6824
rect 95400 6784 95440 6824
rect 3112 6028 3152 6068
rect 3194 6028 3234 6068
rect 3276 6028 3316 6068
rect 3358 6028 3398 6068
rect 3440 6028 3480 6068
rect 18232 6028 18272 6068
rect 18314 6028 18354 6068
rect 18396 6028 18436 6068
rect 18478 6028 18518 6068
rect 18560 6028 18600 6068
rect 33352 6028 33392 6068
rect 33434 6028 33474 6068
rect 33516 6028 33556 6068
rect 33598 6028 33638 6068
rect 33680 6028 33720 6068
rect 48472 6028 48512 6068
rect 48554 6028 48594 6068
rect 48636 6028 48676 6068
rect 48718 6028 48758 6068
rect 48800 6028 48840 6068
rect 63592 6028 63632 6068
rect 63674 6028 63714 6068
rect 63756 6028 63796 6068
rect 63838 6028 63878 6068
rect 63920 6028 63960 6068
rect 78712 6028 78752 6068
rect 78794 6028 78834 6068
rect 78876 6028 78916 6068
rect 78958 6028 78998 6068
rect 79040 6028 79080 6068
rect 93832 6028 93872 6068
rect 93914 6028 93954 6068
rect 93996 6028 94036 6068
rect 94078 6028 94118 6068
rect 94160 6028 94200 6068
rect 844 5692 884 5732
rect 652 5440 692 5480
rect 4352 5272 4392 5312
rect 4434 5272 4474 5312
rect 4516 5272 4556 5312
rect 4598 5272 4638 5312
rect 4680 5272 4720 5312
rect 19472 5272 19512 5312
rect 19554 5272 19594 5312
rect 19636 5272 19676 5312
rect 19718 5272 19758 5312
rect 19800 5272 19840 5312
rect 34592 5272 34632 5312
rect 34674 5272 34714 5312
rect 34756 5272 34796 5312
rect 34838 5272 34878 5312
rect 34920 5272 34960 5312
rect 49712 5272 49752 5312
rect 49794 5272 49834 5312
rect 49876 5272 49916 5312
rect 49958 5272 49998 5312
rect 50040 5272 50080 5312
rect 64832 5272 64872 5312
rect 64914 5272 64954 5312
rect 64996 5272 65036 5312
rect 65078 5272 65118 5312
rect 65160 5272 65200 5312
rect 79952 5272 79992 5312
rect 80034 5272 80074 5312
rect 80116 5272 80156 5312
rect 80198 5272 80238 5312
rect 80280 5272 80320 5312
rect 95072 5272 95112 5312
rect 95154 5272 95194 5312
rect 95236 5272 95276 5312
rect 95318 5272 95358 5312
rect 95400 5272 95440 5312
rect 844 4852 884 4892
rect 652 4768 692 4808
rect 3112 4516 3152 4556
rect 3194 4516 3234 4556
rect 3276 4516 3316 4556
rect 3358 4516 3398 4556
rect 3440 4516 3480 4556
rect 18232 4516 18272 4556
rect 18314 4516 18354 4556
rect 18396 4516 18436 4556
rect 18478 4516 18518 4556
rect 18560 4516 18600 4556
rect 33352 4516 33392 4556
rect 33434 4516 33474 4556
rect 33516 4516 33556 4556
rect 33598 4516 33638 4556
rect 33680 4516 33720 4556
rect 48472 4516 48512 4556
rect 48554 4516 48594 4556
rect 48636 4516 48676 4556
rect 48718 4516 48758 4556
rect 48800 4516 48840 4556
rect 63592 4516 63632 4556
rect 63674 4516 63714 4556
rect 63756 4516 63796 4556
rect 63838 4516 63878 4556
rect 63920 4516 63960 4556
rect 78712 4516 78752 4556
rect 78794 4516 78834 4556
rect 78876 4516 78916 4556
rect 78958 4516 78998 4556
rect 79040 4516 79080 4556
rect 93832 4516 93872 4556
rect 93914 4516 93954 4556
rect 93996 4516 94036 4556
rect 94078 4516 94118 4556
rect 94160 4516 94200 4556
rect 844 4180 884 4220
rect 652 3928 692 3968
rect 4352 3760 4392 3800
rect 4434 3760 4474 3800
rect 4516 3760 4556 3800
rect 4598 3760 4638 3800
rect 4680 3760 4720 3800
rect 19472 3760 19512 3800
rect 19554 3760 19594 3800
rect 19636 3760 19676 3800
rect 19718 3760 19758 3800
rect 19800 3760 19840 3800
rect 34592 3760 34632 3800
rect 34674 3760 34714 3800
rect 34756 3760 34796 3800
rect 34838 3760 34878 3800
rect 34920 3760 34960 3800
rect 49712 3760 49752 3800
rect 49794 3760 49834 3800
rect 49876 3760 49916 3800
rect 49958 3760 49998 3800
rect 50040 3760 50080 3800
rect 64832 3760 64872 3800
rect 64914 3760 64954 3800
rect 64996 3760 65036 3800
rect 65078 3760 65118 3800
rect 65160 3760 65200 3800
rect 79952 3760 79992 3800
rect 80034 3760 80074 3800
rect 80116 3760 80156 3800
rect 80198 3760 80238 3800
rect 80280 3760 80320 3800
rect 95072 3760 95112 3800
rect 95154 3760 95194 3800
rect 95236 3760 95276 3800
rect 95318 3760 95358 3800
rect 95400 3760 95440 3800
rect 844 3340 884 3380
rect 652 3172 692 3212
rect 3112 3004 3152 3044
rect 3194 3004 3234 3044
rect 3276 3004 3316 3044
rect 3358 3004 3398 3044
rect 3440 3004 3480 3044
rect 18232 3004 18272 3044
rect 18314 3004 18354 3044
rect 18396 3004 18436 3044
rect 18478 3004 18518 3044
rect 18560 3004 18600 3044
rect 33352 3004 33392 3044
rect 33434 3004 33474 3044
rect 33516 3004 33556 3044
rect 33598 3004 33638 3044
rect 33680 3004 33720 3044
rect 48472 3004 48512 3044
rect 48554 3004 48594 3044
rect 48636 3004 48676 3044
rect 48718 3004 48758 3044
rect 48800 3004 48840 3044
rect 63592 3004 63632 3044
rect 63674 3004 63714 3044
rect 63756 3004 63796 3044
rect 63838 3004 63878 3044
rect 63920 3004 63960 3044
rect 78712 3004 78752 3044
rect 78794 3004 78834 3044
rect 78876 3004 78916 3044
rect 78958 3004 78998 3044
rect 79040 3004 79080 3044
rect 93832 3004 93872 3044
rect 93914 3004 93954 3044
rect 93996 3004 94036 3044
rect 94078 3004 94118 3044
rect 94160 3004 94200 3044
rect 844 2668 884 2708
rect 652 2416 692 2456
rect 4352 2248 4392 2288
rect 4434 2248 4474 2288
rect 4516 2248 4556 2288
rect 4598 2248 4638 2288
rect 4680 2248 4720 2288
rect 19472 2248 19512 2288
rect 19554 2248 19594 2288
rect 19636 2248 19676 2288
rect 19718 2248 19758 2288
rect 19800 2248 19840 2288
rect 34592 2248 34632 2288
rect 34674 2248 34714 2288
rect 34756 2248 34796 2288
rect 34838 2248 34878 2288
rect 34920 2248 34960 2288
rect 49712 2248 49752 2288
rect 49794 2248 49834 2288
rect 49876 2248 49916 2288
rect 49958 2248 49998 2288
rect 50040 2248 50080 2288
rect 64832 2248 64872 2288
rect 64914 2248 64954 2288
rect 64996 2248 65036 2288
rect 65078 2248 65118 2288
rect 65160 2248 65200 2288
rect 79952 2248 79992 2288
rect 80034 2248 80074 2288
rect 80116 2248 80156 2288
rect 80198 2248 80238 2288
rect 80280 2248 80320 2288
rect 95072 2248 95112 2288
rect 95154 2248 95194 2288
rect 95236 2248 95276 2288
rect 95318 2248 95358 2288
rect 95400 2248 95440 2288
rect 3112 1492 3152 1532
rect 3194 1492 3234 1532
rect 3276 1492 3316 1532
rect 3358 1492 3398 1532
rect 3440 1492 3480 1532
rect 18232 1492 18272 1532
rect 18314 1492 18354 1532
rect 18396 1492 18436 1532
rect 18478 1492 18518 1532
rect 18560 1492 18600 1532
rect 33352 1492 33392 1532
rect 33434 1492 33474 1532
rect 33516 1492 33556 1532
rect 33598 1492 33638 1532
rect 33680 1492 33720 1532
rect 48472 1492 48512 1532
rect 48554 1492 48594 1532
rect 48636 1492 48676 1532
rect 48718 1492 48758 1532
rect 48800 1492 48840 1532
rect 63592 1492 63632 1532
rect 63674 1492 63714 1532
rect 63756 1492 63796 1532
rect 63838 1492 63878 1532
rect 63920 1492 63960 1532
rect 78712 1492 78752 1532
rect 78794 1492 78834 1532
rect 78876 1492 78916 1532
rect 78958 1492 78998 1532
rect 79040 1492 79080 1532
rect 93832 1492 93872 1532
rect 93914 1492 93954 1532
rect 93996 1492 94036 1532
rect 94078 1492 94118 1532
rect 94160 1492 94200 1532
rect 4352 736 4392 776
rect 4434 736 4474 776
rect 4516 736 4556 776
rect 4598 736 4638 776
rect 4680 736 4720 776
rect 19472 736 19512 776
rect 19554 736 19594 776
rect 19636 736 19676 776
rect 19718 736 19758 776
rect 19800 736 19840 776
rect 34592 736 34632 776
rect 34674 736 34714 776
rect 34756 736 34796 776
rect 34838 736 34878 776
rect 34920 736 34960 776
rect 49712 736 49752 776
rect 49794 736 49834 776
rect 49876 736 49916 776
rect 49958 736 49998 776
rect 50040 736 50080 776
rect 64832 736 64872 776
rect 64914 736 64954 776
rect 64996 736 65036 776
rect 65078 736 65118 776
rect 65160 736 65200 776
rect 79952 736 79992 776
rect 80034 736 80074 776
rect 80116 736 80156 776
rect 80198 736 80238 776
rect 80280 736 80320 776
rect 95072 736 95112 776
rect 95154 736 95194 776
rect 95236 736 95276 776
rect 95318 736 95358 776
rect 95400 736 95440 776
<< metal2 >>
rect 4352 38576 4720 38585
rect 4392 38536 4434 38576
rect 4474 38536 4516 38576
rect 4556 38536 4598 38576
rect 4638 38536 4680 38576
rect 4352 38527 4720 38536
rect 19472 38576 19840 38585
rect 19512 38536 19554 38576
rect 19594 38536 19636 38576
rect 19676 38536 19718 38576
rect 19758 38536 19800 38576
rect 19472 38527 19840 38536
rect 34592 38576 34960 38585
rect 34632 38536 34674 38576
rect 34714 38536 34756 38576
rect 34796 38536 34838 38576
rect 34878 38536 34920 38576
rect 34592 38527 34960 38536
rect 49712 38576 50080 38585
rect 49752 38536 49794 38576
rect 49834 38536 49876 38576
rect 49916 38536 49958 38576
rect 49998 38536 50040 38576
rect 49712 38527 50080 38536
rect 64832 38576 65200 38585
rect 64872 38536 64914 38576
rect 64954 38536 64996 38576
rect 65036 38536 65078 38576
rect 65118 38536 65160 38576
rect 64832 38527 65200 38536
rect 79952 38576 80320 38585
rect 79992 38536 80034 38576
rect 80074 38536 80116 38576
rect 80156 38536 80198 38576
rect 80238 38536 80280 38576
rect 79952 38527 80320 38536
rect 95072 38576 95440 38585
rect 95112 38536 95154 38576
rect 95194 38536 95236 38576
rect 95276 38536 95318 38576
rect 95358 38536 95400 38576
rect 95072 38527 95440 38536
rect 3112 37820 3480 37829
rect 3152 37780 3194 37820
rect 3234 37780 3276 37820
rect 3316 37780 3358 37820
rect 3398 37780 3440 37820
rect 3112 37771 3480 37780
rect 18232 37820 18600 37829
rect 18272 37780 18314 37820
rect 18354 37780 18396 37820
rect 18436 37780 18478 37820
rect 18518 37780 18560 37820
rect 18232 37771 18600 37780
rect 33352 37820 33720 37829
rect 33392 37780 33434 37820
rect 33474 37780 33516 37820
rect 33556 37780 33598 37820
rect 33638 37780 33680 37820
rect 33352 37771 33720 37780
rect 48472 37820 48840 37829
rect 48512 37780 48554 37820
rect 48594 37780 48636 37820
rect 48676 37780 48718 37820
rect 48758 37780 48800 37820
rect 48472 37771 48840 37780
rect 63592 37820 63960 37829
rect 63632 37780 63674 37820
rect 63714 37780 63756 37820
rect 63796 37780 63838 37820
rect 63878 37780 63920 37820
rect 63592 37771 63960 37780
rect 78712 37820 79080 37829
rect 78752 37780 78794 37820
rect 78834 37780 78876 37820
rect 78916 37780 78958 37820
rect 78998 37780 79040 37820
rect 78712 37771 79080 37780
rect 93832 37820 94200 37829
rect 93872 37780 93914 37820
rect 93954 37780 93996 37820
rect 94036 37780 94078 37820
rect 94118 37780 94160 37820
rect 93832 37771 94200 37780
rect 267 37568 309 37577
rect 267 37528 268 37568
rect 308 37528 309 37568
rect 267 37519 309 37528
rect 75 36728 117 36737
rect 75 36688 76 36728
rect 116 36688 117 36728
rect 75 36679 117 36688
rect 76 32780 116 36679
rect 76 32740 212 32780
rect 172 21617 212 32740
rect 268 26237 308 37519
rect 4352 37064 4720 37073
rect 4392 37024 4434 37064
rect 4474 37024 4516 37064
rect 4556 37024 4598 37064
rect 4638 37024 4680 37064
rect 4352 37015 4720 37024
rect 19472 37064 19840 37073
rect 19512 37024 19554 37064
rect 19594 37024 19636 37064
rect 19676 37024 19718 37064
rect 19758 37024 19800 37064
rect 19472 37015 19840 37024
rect 34592 37064 34960 37073
rect 34632 37024 34674 37064
rect 34714 37024 34756 37064
rect 34796 37024 34838 37064
rect 34878 37024 34920 37064
rect 34592 37015 34960 37024
rect 49712 37064 50080 37073
rect 49752 37024 49794 37064
rect 49834 37024 49876 37064
rect 49916 37024 49958 37064
rect 49998 37024 50040 37064
rect 49712 37015 50080 37024
rect 64832 37064 65200 37073
rect 64872 37024 64914 37064
rect 64954 37024 64996 37064
rect 65036 37024 65078 37064
rect 65118 37024 65160 37064
rect 64832 37015 65200 37024
rect 79952 37064 80320 37073
rect 79992 37024 80034 37064
rect 80074 37024 80116 37064
rect 80156 37024 80198 37064
rect 80238 37024 80280 37064
rect 79952 37015 80320 37024
rect 95072 37064 95440 37073
rect 95112 37024 95154 37064
rect 95194 37024 95236 37064
rect 95276 37024 95318 37064
rect 95358 37024 95400 37064
rect 95072 37015 95440 37024
rect 3112 36308 3480 36317
rect 3152 36268 3194 36308
rect 3234 36268 3276 36308
rect 3316 36268 3358 36308
rect 3398 36268 3440 36308
rect 3112 36259 3480 36268
rect 18232 36308 18600 36317
rect 18272 36268 18314 36308
rect 18354 36268 18396 36308
rect 18436 36268 18478 36308
rect 18518 36268 18560 36308
rect 18232 36259 18600 36268
rect 33352 36308 33720 36317
rect 33392 36268 33434 36308
rect 33474 36268 33516 36308
rect 33556 36268 33598 36308
rect 33638 36268 33680 36308
rect 33352 36259 33720 36268
rect 48472 36308 48840 36317
rect 48512 36268 48554 36308
rect 48594 36268 48636 36308
rect 48676 36268 48718 36308
rect 48758 36268 48800 36308
rect 48472 36259 48840 36268
rect 63592 36308 63960 36317
rect 63632 36268 63674 36308
rect 63714 36268 63756 36308
rect 63796 36268 63838 36308
rect 63878 36268 63920 36308
rect 63592 36259 63960 36268
rect 78712 36308 79080 36317
rect 78752 36268 78794 36308
rect 78834 36268 78876 36308
rect 78916 36268 78958 36308
rect 78998 36268 79040 36308
rect 78712 36259 79080 36268
rect 93832 36308 94200 36317
rect 93872 36268 93914 36308
rect 93954 36268 93996 36308
rect 94036 36268 94078 36308
rect 94118 36268 94160 36308
rect 93832 36259 94200 36268
rect 4352 35552 4720 35561
rect 4392 35512 4434 35552
rect 4474 35512 4516 35552
rect 4556 35512 4598 35552
rect 4638 35512 4680 35552
rect 4352 35503 4720 35512
rect 19472 35552 19840 35561
rect 19512 35512 19554 35552
rect 19594 35512 19636 35552
rect 19676 35512 19718 35552
rect 19758 35512 19800 35552
rect 19472 35503 19840 35512
rect 34592 35552 34960 35561
rect 34632 35512 34674 35552
rect 34714 35512 34756 35552
rect 34796 35512 34838 35552
rect 34878 35512 34920 35552
rect 34592 35503 34960 35512
rect 49712 35552 50080 35561
rect 49752 35512 49794 35552
rect 49834 35512 49876 35552
rect 49916 35512 49958 35552
rect 49998 35512 50040 35552
rect 49712 35503 50080 35512
rect 64832 35552 65200 35561
rect 64872 35512 64914 35552
rect 64954 35512 64996 35552
rect 65036 35512 65078 35552
rect 65118 35512 65160 35552
rect 64832 35503 65200 35512
rect 79952 35552 80320 35561
rect 79992 35512 80034 35552
rect 80074 35512 80116 35552
rect 80156 35512 80198 35552
rect 80238 35512 80280 35552
rect 79952 35503 80320 35512
rect 95072 35552 95440 35561
rect 95112 35512 95154 35552
rect 95194 35512 95236 35552
rect 95276 35512 95318 35552
rect 95358 35512 95400 35552
rect 95072 35503 95440 35512
rect 652 35216 692 35225
rect 652 35057 692 35176
rect 843 35216 885 35225
rect 843 35176 844 35216
rect 884 35176 885 35216
rect 843 35167 885 35176
rect 23499 35216 23541 35225
rect 23499 35176 23500 35216
rect 23540 35176 23541 35216
rect 23499 35167 23541 35176
rect 844 35082 884 35167
rect 651 35048 693 35057
rect 651 35008 652 35048
rect 692 35008 693 35048
rect 651 34999 693 35008
rect 3112 34796 3480 34805
rect 3152 34756 3194 34796
rect 3234 34756 3276 34796
rect 3316 34756 3358 34796
rect 3398 34756 3440 34796
rect 3112 34747 3480 34756
rect 18232 34796 18600 34805
rect 18272 34756 18314 34796
rect 18354 34756 18396 34796
rect 18436 34756 18478 34796
rect 18518 34756 18560 34796
rect 18232 34747 18600 34756
rect 652 34376 692 34385
rect 652 34217 692 34336
rect 843 34376 885 34385
rect 843 34336 844 34376
rect 884 34336 885 34376
rect 843 34327 885 34336
rect 844 34242 884 34327
rect 651 34208 693 34217
rect 651 34168 652 34208
rect 692 34168 693 34208
rect 651 34159 693 34168
rect 4352 34040 4720 34049
rect 4392 34000 4434 34040
rect 4474 34000 4516 34040
rect 4556 34000 4598 34040
rect 4638 34000 4680 34040
rect 4352 33991 4720 34000
rect 19472 34040 19840 34049
rect 19512 34000 19554 34040
rect 19594 34000 19636 34040
rect 19676 34000 19718 34040
rect 19758 34000 19800 34040
rect 19472 33991 19840 34000
rect 652 33704 692 33713
rect 652 33377 692 33664
rect 843 33704 885 33713
rect 843 33664 844 33704
rect 884 33664 885 33704
rect 843 33655 885 33664
rect 844 33570 884 33655
rect 651 33368 693 33377
rect 651 33328 652 33368
rect 692 33328 693 33368
rect 651 33319 693 33328
rect 3112 33284 3480 33293
rect 3152 33244 3194 33284
rect 3234 33244 3276 33284
rect 3316 33244 3358 33284
rect 3398 33244 3440 33284
rect 3112 33235 3480 33244
rect 18232 33284 18600 33293
rect 18272 33244 18314 33284
rect 18354 33244 18396 33284
rect 18436 33244 18478 33284
rect 18518 33244 18560 33284
rect 18232 33235 18600 33244
rect 844 32873 884 32958
rect 652 32864 692 32873
rect 652 32537 692 32824
rect 843 32864 885 32873
rect 843 32824 844 32864
rect 884 32824 885 32864
rect 843 32815 885 32824
rect 651 32528 693 32537
rect 651 32488 652 32528
rect 692 32488 693 32528
rect 651 32479 693 32488
rect 4352 32528 4720 32537
rect 4392 32488 4434 32528
rect 4474 32488 4516 32528
rect 4556 32488 4598 32528
rect 4638 32488 4680 32528
rect 4352 32479 4720 32488
rect 19472 32528 19840 32537
rect 19512 32488 19554 32528
rect 19594 32488 19636 32528
rect 19676 32488 19718 32528
rect 19758 32488 19800 32528
rect 19472 32479 19840 32488
rect 652 32108 692 32117
rect 652 31697 692 32068
rect 844 31940 884 31949
rect 884 31900 1172 31940
rect 844 31891 884 31900
rect 651 31688 693 31697
rect 651 31648 652 31688
rect 692 31648 693 31688
rect 651 31639 693 31648
rect 652 31436 692 31445
rect 652 30857 692 31396
rect 844 31184 884 31193
rect 884 31144 1076 31184
rect 844 31135 884 31144
rect 651 30848 693 30857
rect 651 30808 652 30848
rect 692 30808 693 30848
rect 651 30799 693 30808
rect 652 30596 692 30605
rect 652 30101 692 30556
rect 844 30428 884 30437
rect 748 30388 844 30428
rect 651 30092 693 30101
rect 651 30052 652 30092
rect 692 30052 693 30092
rect 651 30043 693 30052
rect 652 29924 692 29933
rect 652 29177 692 29884
rect 651 29168 693 29177
rect 651 29128 652 29168
rect 692 29128 693 29168
rect 651 29119 693 29128
rect 651 28328 693 28337
rect 651 28288 652 28328
rect 692 28288 693 28328
rect 651 28279 693 28288
rect 652 28194 692 28279
rect 748 27833 788 30388
rect 844 30379 884 30388
rect 844 29672 884 29681
rect 884 29632 980 29672
rect 844 29623 884 29632
rect 843 28328 885 28337
rect 843 28288 844 28328
rect 884 28288 885 28328
rect 843 28279 885 28288
rect 844 28194 884 28279
rect 747 27824 789 27833
rect 747 27784 748 27824
rect 788 27784 789 27824
rect 747 27775 789 27784
rect 652 27656 692 27665
rect 652 27497 692 27616
rect 844 27656 884 27665
rect 651 27488 693 27497
rect 651 27448 652 27488
rect 692 27448 693 27488
rect 651 27439 693 27448
rect 844 26984 884 27616
rect 940 27497 980 29632
rect 939 27488 981 27497
rect 939 27448 940 27488
rect 980 27448 981 27488
rect 939 27439 981 27448
rect 1036 26993 1076 31144
rect 1132 29849 1172 31900
rect 3112 31772 3480 31781
rect 3152 31732 3194 31772
rect 3234 31732 3276 31772
rect 3316 31732 3358 31772
rect 3398 31732 3440 31772
rect 3112 31723 3480 31732
rect 18232 31772 18600 31781
rect 18272 31732 18314 31772
rect 18354 31732 18396 31772
rect 18436 31732 18478 31772
rect 18518 31732 18560 31772
rect 18232 31723 18600 31732
rect 21772 31352 21812 31361
rect 21772 31277 21812 31312
rect 22635 31352 22677 31361
rect 22635 31312 22636 31352
rect 22676 31312 22677 31352
rect 22635 31303 22677 31312
rect 21388 31268 21428 31277
rect 4352 31016 4720 31025
rect 4392 30976 4434 31016
rect 4474 30976 4516 31016
rect 4556 30976 4598 31016
rect 4638 30976 4680 31016
rect 4352 30967 4720 30976
rect 19472 31016 19840 31025
rect 19512 30976 19554 31016
rect 19594 30976 19636 31016
rect 19676 30976 19718 31016
rect 19758 30976 19800 31016
rect 19472 30967 19840 30976
rect 3112 30260 3480 30269
rect 3152 30220 3194 30260
rect 3234 30220 3276 30260
rect 3316 30220 3358 30260
rect 3398 30220 3440 30260
rect 3112 30211 3480 30220
rect 18232 30260 18600 30269
rect 18272 30220 18314 30260
rect 18354 30220 18396 30260
rect 18436 30220 18478 30260
rect 18518 30220 18560 30260
rect 18232 30211 18600 30220
rect 1131 29840 1173 29849
rect 1131 29800 1132 29840
rect 1172 29800 1173 29840
rect 1131 29791 1173 29800
rect 19947 29840 19989 29849
rect 19947 29800 19948 29840
rect 19988 29800 19989 29840
rect 19947 29791 19989 29800
rect 4352 29504 4720 29513
rect 4392 29464 4434 29504
rect 4474 29464 4516 29504
rect 4556 29464 4598 29504
rect 4638 29464 4680 29504
rect 4352 29455 4720 29464
rect 19472 29504 19840 29513
rect 19512 29464 19554 29504
rect 19594 29464 19636 29504
rect 19676 29464 19718 29504
rect 19758 29464 19800 29504
rect 19472 29455 19840 29464
rect 15340 29168 15380 29177
rect 15724 29168 15764 29177
rect 3112 28748 3480 28757
rect 3152 28708 3194 28748
rect 3234 28708 3276 28748
rect 3316 28708 3358 28748
rect 3398 28708 3440 28748
rect 3112 28699 3480 28708
rect 15340 28337 15380 29128
rect 15436 29128 15724 29168
rect 15339 28328 15381 28337
rect 15339 28288 15340 28328
rect 15380 28288 15381 28328
rect 15339 28279 15381 28288
rect 4352 27992 4720 28001
rect 4392 27952 4434 27992
rect 4474 27952 4516 27992
rect 4556 27952 4598 27992
rect 4638 27952 4680 27992
rect 4352 27943 4720 27952
rect 3112 27236 3480 27245
rect 3152 27196 3194 27236
rect 3234 27196 3276 27236
rect 3316 27196 3358 27236
rect 3398 27196 3440 27236
rect 3112 27187 3480 27196
rect 1035 26984 1077 26993
rect 844 26944 980 26984
rect 652 26816 692 26825
rect 844 26816 884 26825
rect 652 26657 692 26776
rect 748 26776 844 26816
rect 651 26648 693 26657
rect 651 26608 652 26648
rect 692 26608 693 26648
rect 651 26599 693 26608
rect 748 26312 788 26776
rect 844 26767 884 26776
rect 556 26272 788 26312
rect 267 26228 309 26237
rect 267 26188 268 26228
rect 308 26188 309 26228
rect 267 26179 309 26188
rect 171 21608 213 21617
rect 171 21568 172 21608
rect 212 21568 213 21608
rect 171 21559 213 21568
rect 556 19853 596 26272
rect 652 26144 692 26153
rect 844 26144 884 26153
rect 652 25817 692 26104
rect 748 26104 844 26144
rect 651 25808 693 25817
rect 651 25768 652 25808
rect 692 25768 693 25808
rect 651 25759 693 25768
rect 652 25304 692 25313
rect 652 24977 692 25264
rect 651 24968 693 24977
rect 651 24928 652 24968
rect 692 24928 693 24968
rect 651 24919 693 24928
rect 652 24632 692 24641
rect 652 24137 692 24592
rect 651 24128 693 24137
rect 651 24088 652 24128
rect 692 24088 693 24128
rect 651 24079 693 24088
rect 652 23792 692 23801
rect 652 23297 692 23752
rect 651 23288 693 23297
rect 651 23248 652 23288
rect 692 23248 693 23288
rect 651 23239 693 23248
rect 652 22448 692 22457
rect 652 21701 692 22408
rect 651 21692 693 21701
rect 651 21652 652 21692
rect 692 21652 693 21692
rect 651 21643 693 21652
rect 652 20936 692 20945
rect 652 20777 692 20896
rect 651 20768 693 20777
rect 651 20728 652 20768
rect 692 20728 693 20768
rect 651 20719 693 20728
rect 748 20021 788 26104
rect 844 26095 884 26104
rect 940 25481 980 26944
rect 1035 26944 1036 26984
rect 1076 26944 1077 26984
rect 1035 26935 1077 26944
rect 14859 26648 14901 26657
rect 14859 26608 14860 26648
rect 14900 26608 14901 26648
rect 14859 26599 14901 26608
rect 4352 26480 4720 26489
rect 4392 26440 4434 26480
rect 4474 26440 4516 26480
rect 4556 26440 4598 26480
rect 4638 26440 4680 26480
rect 4352 26431 4720 26440
rect 14860 26228 14900 26599
rect 14860 26179 14900 26188
rect 15244 26144 15284 26153
rect 15436 26144 15476 29128
rect 15724 29119 15764 29128
rect 16588 29168 16628 29177
rect 16588 26405 16628 29128
rect 17740 28916 17780 28925
rect 17780 28876 18164 28916
rect 17740 28867 17780 28876
rect 18124 28244 18164 28876
rect 18232 28748 18600 28757
rect 18272 28708 18314 28748
rect 18354 28708 18396 28748
rect 18436 28708 18478 28748
rect 18518 28708 18560 28748
rect 18232 28699 18600 28708
rect 18124 28204 18452 28244
rect 18219 28076 18261 28085
rect 18219 28036 18220 28076
rect 18260 28036 18261 28076
rect 18219 28027 18261 28036
rect 17259 27656 17301 27665
rect 17259 27616 17260 27656
rect 17300 27616 17301 27656
rect 17259 27607 17301 27616
rect 18123 27656 18165 27665
rect 18123 27616 18124 27656
rect 18164 27616 18165 27656
rect 18123 27607 18165 27616
rect 16107 26396 16149 26405
rect 16107 26356 16108 26396
rect 16148 26356 16149 26396
rect 16107 26347 16149 26356
rect 16587 26396 16629 26405
rect 16587 26356 16588 26396
rect 16628 26356 16629 26396
rect 16587 26347 16629 26356
rect 15284 26104 15476 26144
rect 16108 26144 16148 26347
rect 17260 26312 17300 27607
rect 18124 27522 18164 27607
rect 18220 27572 18260 28027
rect 18220 27523 18260 27532
rect 18412 27572 18452 28204
rect 19472 27992 19840 28001
rect 19512 27952 19554 27992
rect 19594 27952 19636 27992
rect 19676 27952 19718 27992
rect 19758 27952 19800 27992
rect 19472 27943 19840 27952
rect 19948 27824 19988 29791
rect 21388 28589 21428 31228
rect 21771 31268 21813 31277
rect 21771 31228 21772 31268
rect 21812 31228 21813 31268
rect 21771 31219 21813 31228
rect 21772 28832 21812 31219
rect 21772 28792 21908 28832
rect 21387 28580 21429 28589
rect 21387 28540 21388 28580
rect 21428 28540 21429 28580
rect 21387 28531 21429 28540
rect 19852 27784 19988 27824
rect 20043 27824 20085 27833
rect 20043 27784 20044 27824
rect 20084 27784 20085 27824
rect 18507 27656 18549 27665
rect 18507 27616 18508 27656
rect 18548 27616 18549 27656
rect 18507 27607 18549 27616
rect 18700 27656 18740 27665
rect 18412 27523 18452 27532
rect 18508 27522 18548 27607
rect 18316 27488 18356 27497
rect 18316 27404 18356 27448
rect 18700 27404 18740 27616
rect 18316 27364 18740 27404
rect 18796 27404 18836 27413
rect 18232 27236 18600 27245
rect 18272 27196 18314 27236
rect 18354 27196 18396 27236
rect 18436 27196 18478 27236
rect 18518 27196 18560 27236
rect 18232 27187 18600 27196
rect 17260 26263 17300 26272
rect 3112 25724 3480 25733
rect 3152 25684 3194 25724
rect 3234 25684 3276 25724
rect 3316 25684 3358 25724
rect 3398 25684 3440 25724
rect 3112 25675 3480 25684
rect 939 25472 981 25481
rect 939 25432 940 25472
rect 980 25432 981 25472
rect 939 25423 981 25432
rect 844 25304 884 25313
rect 884 25264 1076 25304
rect 844 25255 884 25264
rect 844 24632 884 24641
rect 844 23960 884 24592
rect 844 23920 980 23960
rect 843 23792 885 23801
rect 843 23752 844 23792
rect 884 23752 885 23792
rect 843 23743 885 23752
rect 844 23658 884 23743
rect 940 20777 980 23920
rect 939 20768 981 20777
rect 939 20728 940 20768
rect 980 20728 981 20768
rect 939 20719 981 20728
rect 747 20012 789 20021
rect 747 19972 748 20012
rect 788 19972 789 20012
rect 747 19963 789 19972
rect 651 19928 693 19937
rect 651 19888 652 19928
rect 692 19888 693 19928
rect 651 19879 693 19888
rect 555 19844 597 19853
rect 555 19804 556 19844
rect 596 19804 597 19844
rect 555 19795 597 19804
rect 652 19794 692 19879
rect 1036 19517 1076 25264
rect 4352 24968 4720 24977
rect 4392 24928 4434 24968
rect 4474 24928 4516 24968
rect 4556 24928 4598 24968
rect 4638 24928 4680 24968
rect 4352 24919 4720 24928
rect 3112 24212 3480 24221
rect 3152 24172 3194 24212
rect 3234 24172 3276 24212
rect 3316 24172 3358 24212
rect 3398 24172 3440 24212
rect 3112 24163 3480 24172
rect 4352 23456 4720 23465
rect 4392 23416 4434 23456
rect 4474 23416 4516 23456
rect 4556 23416 4598 23456
rect 4638 23416 4680 23456
rect 4352 23407 4720 23416
rect 15244 23129 15284 26104
rect 16108 23960 16148 26104
rect 18232 25724 18600 25733
rect 18272 25684 18314 25724
rect 18354 25684 18396 25724
rect 18436 25684 18478 25724
rect 18518 25684 18560 25724
rect 18232 25675 18600 25684
rect 18232 24212 18600 24221
rect 18272 24172 18314 24212
rect 18354 24172 18396 24212
rect 18436 24172 18478 24212
rect 18518 24172 18560 24212
rect 18232 24163 18600 24172
rect 18796 23960 18836 27364
rect 19852 26816 19892 27784
rect 20043 27775 20085 27784
rect 21483 27824 21525 27833
rect 21483 27784 21484 27824
rect 21524 27784 21525 27824
rect 21483 27775 21525 27784
rect 20044 27690 20084 27775
rect 20140 27656 20180 27665
rect 20140 27497 20180 27616
rect 20235 27656 20277 27665
rect 20235 27616 20236 27656
rect 20276 27616 20277 27656
rect 20235 27607 20277 27616
rect 20139 27488 20181 27497
rect 20139 27448 20140 27488
rect 20180 27448 20181 27488
rect 20139 27439 20181 27448
rect 19948 26993 19988 27078
rect 19947 26984 19989 26993
rect 19947 26944 19948 26984
rect 19988 26944 19989 26984
rect 19947 26935 19989 26944
rect 20236 26909 20276 27607
rect 20332 27404 20372 27413
rect 20372 27364 20564 27404
rect 20332 27355 20372 27364
rect 20428 26909 20468 26911
rect 20235 26900 20277 26909
rect 20235 26860 20236 26900
rect 20276 26860 20277 26900
rect 20235 26851 20277 26860
rect 20427 26900 20469 26909
rect 20427 26860 20428 26900
rect 20468 26860 20469 26900
rect 20427 26851 20469 26860
rect 19948 26816 19988 26825
rect 19852 26776 19948 26816
rect 19948 26767 19988 26776
rect 20139 26816 20181 26825
rect 20139 26776 20140 26816
rect 20180 26776 20181 26816
rect 20139 26767 20181 26776
rect 20428 26816 20468 26851
rect 20428 26767 20468 26776
rect 20524 26816 20564 27364
rect 20524 26767 20564 26776
rect 20619 26816 20661 26825
rect 20619 26776 20620 26816
rect 20660 26776 20661 26816
rect 20619 26767 20661 26776
rect 20140 26648 20180 26767
rect 20620 26682 20660 26767
rect 20140 26599 20180 26608
rect 20331 26648 20373 26657
rect 20331 26608 20332 26648
rect 20372 26608 20373 26648
rect 20331 26599 20373 26608
rect 20332 26514 20372 26599
rect 19472 26480 19840 26489
rect 19512 26440 19554 26480
rect 19594 26440 19636 26480
rect 19676 26440 19718 26480
rect 19758 26440 19800 26480
rect 19472 26431 19840 26440
rect 21484 26144 21524 27775
rect 21579 27740 21621 27749
rect 21579 27700 21580 27740
rect 21620 27700 21621 27740
rect 21579 27691 21621 27700
rect 21580 26312 21620 27691
rect 21675 27488 21717 27497
rect 21675 27448 21676 27488
rect 21716 27448 21717 27488
rect 21675 27439 21717 27448
rect 21580 26263 21620 26272
rect 21484 26095 21524 26104
rect 21676 26144 21716 27439
rect 21771 26816 21813 26825
rect 21771 26776 21772 26816
rect 21812 26776 21813 26816
rect 21771 26767 21813 26776
rect 21676 26095 21716 26104
rect 21772 26144 21812 26767
rect 21772 26095 21812 26104
rect 19472 24968 19840 24977
rect 19512 24928 19554 24968
rect 19594 24928 19636 24968
rect 19676 24928 19718 24968
rect 19758 24928 19800 24968
rect 19472 24919 19840 24928
rect 16108 23920 16244 23960
rect 15243 23120 15285 23129
rect 15243 23080 15244 23120
rect 15284 23080 15285 23120
rect 15243 23071 15285 23080
rect 3112 22700 3480 22709
rect 3152 22660 3194 22700
rect 3234 22660 3276 22700
rect 3316 22660 3358 22700
rect 3398 22660 3440 22700
rect 3112 22651 3480 22660
rect 15244 22280 15284 23071
rect 15340 22280 15380 22289
rect 15244 22240 15340 22280
rect 15340 22231 15380 22240
rect 16204 22280 16244 23920
rect 16204 22231 16244 22240
rect 18124 23920 18836 23960
rect 14956 22196 14996 22205
rect 4352 21944 4720 21953
rect 4392 21904 4434 21944
rect 4474 21904 4516 21944
rect 4556 21904 4598 21944
rect 4638 21904 4680 21944
rect 4352 21895 4720 21904
rect 3112 21188 3480 21197
rect 3152 21148 3194 21188
rect 3234 21148 3276 21188
rect 3316 21148 3358 21188
rect 3398 21148 3440 21188
rect 3112 21139 3480 21148
rect 1131 20516 1173 20525
rect 1131 20476 1132 20516
rect 1172 20476 1173 20516
rect 1131 20467 1173 20476
rect 1035 19508 1077 19517
rect 1035 19468 1036 19508
rect 1076 19468 1077 19508
rect 1035 19459 1077 19468
rect 652 19424 692 19433
rect 652 19097 692 19384
rect 651 19088 693 19097
rect 651 19048 652 19088
rect 692 19048 693 19088
rect 651 19039 693 19048
rect 652 18416 692 18425
rect 652 18257 692 18376
rect 651 18248 693 18257
rect 651 18208 652 18248
rect 692 18208 693 18248
rect 651 18199 693 18208
rect 652 17912 692 17921
rect 652 17417 692 17872
rect 651 17408 693 17417
rect 651 17368 652 17408
rect 692 17368 693 17408
rect 651 17359 693 17368
rect 652 16904 692 16913
rect 652 16577 692 16864
rect 651 16568 693 16577
rect 651 16528 652 16568
rect 692 16528 693 16568
rect 651 16519 693 16528
rect 652 16400 692 16409
rect 556 16360 652 16400
rect 556 15737 596 16360
rect 652 16351 692 16360
rect 555 15728 597 15737
rect 555 15688 556 15728
rect 596 15688 597 15728
rect 555 15679 597 15688
rect 652 15728 692 15737
rect 652 14897 692 15688
rect 939 15308 981 15317
rect 939 15268 940 15308
rect 980 15268 981 15308
rect 939 15259 981 15268
rect 651 14888 693 14897
rect 651 14848 652 14888
rect 692 14848 693 14888
rect 651 14839 693 14848
rect 652 14552 692 14561
rect 652 14057 692 14512
rect 651 14048 693 14057
rect 651 14008 652 14048
rect 692 14008 693 14048
rect 651 13999 693 14008
rect 651 13208 693 13217
rect 651 13168 652 13208
rect 692 13168 693 13208
rect 651 13159 693 13168
rect 652 13040 692 13159
rect 652 12991 692 13000
rect 843 13040 885 13049
rect 843 13000 844 13040
rect 884 13000 885 13040
rect 843 12991 885 13000
rect 652 12704 692 12713
rect 652 12377 692 12664
rect 651 12368 693 12377
rect 651 12328 652 12368
rect 692 12328 693 12368
rect 651 12319 693 12328
rect 747 12200 789 12209
rect 747 12160 748 12200
rect 788 12160 789 12200
rect 747 12151 789 12160
rect 651 11528 693 11537
rect 651 11488 652 11528
rect 692 11488 693 11528
rect 651 11479 693 11488
rect 652 11394 692 11479
rect 651 10772 693 10781
rect 651 10732 652 10772
rect 692 10732 693 10772
rect 651 10723 693 10732
rect 652 10638 692 10723
rect 652 10016 692 10025
rect 652 9857 692 9976
rect 651 9848 693 9857
rect 651 9808 652 9848
rect 692 9808 693 9848
rect 651 9799 693 9808
rect 652 9260 692 9269
rect 652 9017 692 9220
rect 651 9008 693 9017
rect 651 8968 652 9008
rect 692 8968 693 9008
rect 651 8959 693 8968
rect 748 8756 788 12151
rect 844 11780 884 12991
rect 844 11731 884 11740
rect 843 10940 885 10949
rect 843 10900 844 10940
rect 884 10900 885 10940
rect 843 10891 885 10900
rect 844 10806 884 10891
rect 843 10268 885 10277
rect 843 10228 844 10268
rect 884 10228 885 10268
rect 843 10219 885 10228
rect 844 10134 884 10219
rect 843 9428 885 9437
rect 843 9388 844 9428
rect 884 9388 885 9428
rect 843 9379 885 9388
rect 844 9294 884 9379
rect 844 8756 884 8765
rect 748 8716 844 8756
rect 844 8707 884 8716
rect 940 8588 980 15259
rect 1035 12032 1077 12041
rect 1035 11992 1036 12032
rect 1076 11992 1077 12032
rect 1035 11983 1077 11992
rect 748 8548 980 8588
rect 652 8504 692 8513
rect 652 8177 692 8464
rect 651 8168 693 8177
rect 651 8128 652 8168
rect 692 8128 693 8168
rect 651 8119 693 8128
rect 652 7748 692 7757
rect 652 7337 692 7708
rect 651 7328 693 7337
rect 651 7288 652 7328
rect 692 7288 693 7328
rect 651 7279 693 7288
rect 652 6992 692 7001
rect 652 6497 692 6952
rect 651 6488 693 6497
rect 651 6448 652 6488
rect 692 6448 693 6488
rect 651 6439 693 6448
rect 651 5648 693 5657
rect 651 5608 652 5648
rect 692 5608 693 5648
rect 651 5599 693 5608
rect 652 5480 692 5599
rect 652 5431 692 5440
rect 651 4808 693 4817
rect 651 4768 652 4808
rect 692 4768 693 4808
rect 651 4759 693 4768
rect 652 4674 692 4759
rect 651 3968 693 3977
rect 651 3928 652 3968
rect 692 3928 693 3968
rect 651 3919 693 3928
rect 652 3834 692 3919
rect 651 3212 693 3221
rect 651 3172 652 3212
rect 692 3172 693 3212
rect 651 3163 693 3172
rect 652 3078 692 3163
rect 748 2708 788 8548
rect 844 7916 884 7925
rect 1036 7916 1076 11983
rect 884 7876 1076 7916
rect 844 7867 884 7876
rect 843 7244 885 7253
rect 843 7204 844 7244
rect 884 7204 885 7244
rect 843 7195 885 7204
rect 844 7110 884 7195
rect 843 5732 885 5741
rect 843 5692 844 5732
rect 884 5692 885 5732
rect 843 5683 885 5692
rect 844 5598 884 5683
rect 843 4892 885 4901
rect 843 4852 844 4892
rect 884 4852 885 4892
rect 843 4843 885 4852
rect 844 4758 884 4843
rect 843 4220 885 4229
rect 843 4180 844 4220
rect 884 4180 885 4220
rect 843 4171 885 4180
rect 844 4086 884 4171
rect 844 3380 884 3389
rect 1132 3380 1172 20467
rect 4352 20432 4720 20441
rect 4392 20392 4434 20432
rect 4474 20392 4516 20432
rect 4556 20392 4598 20432
rect 4638 20392 4680 20432
rect 4352 20383 4720 20392
rect 14956 20189 14996 22156
rect 17355 22112 17397 22121
rect 17355 22072 17356 22112
rect 17396 22072 17397 22112
rect 17355 22063 17397 22072
rect 17356 21978 17396 22063
rect 17739 20768 17781 20777
rect 17739 20728 17740 20768
rect 17780 20728 17781 20768
rect 17739 20719 17781 20728
rect 14955 20180 14997 20189
rect 14955 20140 14956 20180
rect 14996 20140 14997 20180
rect 14955 20131 14997 20140
rect 15435 20180 15477 20189
rect 15435 20140 15436 20180
rect 15476 20140 15477 20180
rect 15435 20131 15477 20140
rect 15436 20046 15476 20131
rect 15628 20096 15668 20105
rect 15628 19937 15668 20056
rect 15916 20096 15956 20105
rect 15916 20021 15956 20056
rect 15915 20012 15957 20021
rect 15915 19972 15916 20012
rect 15956 19972 15957 20012
rect 15915 19963 15957 19972
rect 15627 19928 15669 19937
rect 15627 19888 15628 19928
rect 15668 19888 15669 19928
rect 15627 19879 15669 19888
rect 3112 19676 3480 19685
rect 3152 19636 3194 19676
rect 3234 19636 3276 19676
rect 3316 19636 3358 19676
rect 3398 19636 3440 19676
rect 3112 19627 3480 19636
rect 15628 19172 15668 19879
rect 15916 19265 15956 19963
rect 15915 19256 15957 19265
rect 15915 19216 15916 19256
rect 15956 19216 15957 19256
rect 15915 19207 15957 19216
rect 16107 19256 16149 19265
rect 16107 19216 16108 19256
rect 16148 19216 16149 19256
rect 16107 19207 16149 19216
rect 15723 19172 15765 19181
rect 15628 19132 15724 19172
rect 15764 19132 15765 19172
rect 15723 19123 15765 19132
rect 4352 18920 4720 18929
rect 4392 18880 4434 18920
rect 4474 18880 4516 18920
rect 4556 18880 4598 18920
rect 4638 18880 4680 18920
rect 4352 18871 4720 18880
rect 3112 18164 3480 18173
rect 3152 18124 3194 18164
rect 3234 18124 3276 18164
rect 3316 18124 3358 18164
rect 3398 18124 3440 18164
rect 3112 18115 3480 18124
rect 4352 17408 4720 17417
rect 4392 17368 4434 17408
rect 4474 17368 4516 17408
rect 4556 17368 4598 17408
rect 4638 17368 4680 17408
rect 4352 17359 4720 17368
rect 15724 17072 15764 19123
rect 16108 17744 16148 19207
rect 17548 18668 17588 18677
rect 17588 18628 17684 18668
rect 17548 18619 17588 18628
rect 17644 17753 17684 18628
rect 17740 18584 17780 20719
rect 18027 19508 18069 19517
rect 18027 19468 18028 19508
rect 18068 19468 18069 19508
rect 18027 19459 18069 19468
rect 17740 18535 17780 18544
rect 18028 18584 18068 19459
rect 18028 18535 18068 18544
rect 16108 17695 16148 17704
rect 16203 17744 16245 17753
rect 16203 17704 16204 17744
rect 16244 17704 16245 17744
rect 16203 17695 16245 17704
rect 17643 17744 17685 17753
rect 17643 17704 17644 17744
rect 17684 17704 17685 17744
rect 17643 17695 17685 17704
rect 16204 17610 16244 17695
rect 15820 17576 15860 17585
rect 15860 17536 16052 17576
rect 15820 17527 15860 17536
rect 15820 17072 15860 17081
rect 15724 17032 15820 17072
rect 15820 17023 15860 17032
rect 16012 17072 16052 17536
rect 16012 17023 16052 17032
rect 15916 16988 15956 16997
rect 3112 16652 3480 16661
rect 3152 16612 3194 16652
rect 3234 16612 3276 16652
rect 3316 16612 3358 16652
rect 3398 16612 3440 16652
rect 3112 16603 3480 16612
rect 15916 16232 15956 16948
rect 15436 16192 15956 16232
rect 4352 15896 4720 15905
rect 4392 15856 4434 15896
rect 4474 15856 4516 15896
rect 4556 15856 4598 15896
rect 4638 15856 4680 15896
rect 4352 15847 4720 15856
rect 15436 15644 15476 16192
rect 15436 15595 15476 15604
rect 15820 15560 15860 15569
rect 3112 15140 3480 15149
rect 3152 15100 3194 15140
rect 3234 15100 3276 15140
rect 3316 15100 3358 15140
rect 3398 15100 3440 15140
rect 3112 15091 3480 15100
rect 4352 14384 4720 14393
rect 4392 14344 4434 14384
rect 4474 14344 4516 14384
rect 4556 14344 4598 14384
rect 4638 14344 4680 14384
rect 4352 14335 4720 14344
rect 3112 13628 3480 13637
rect 3152 13588 3194 13628
rect 3234 13588 3276 13628
rect 3316 13588 3358 13628
rect 3398 13588 3440 13628
rect 3112 13579 3480 13588
rect 4352 12872 4720 12881
rect 4392 12832 4434 12872
rect 4474 12832 4516 12872
rect 4556 12832 4598 12872
rect 4638 12832 4680 12872
rect 4352 12823 4720 12832
rect 15820 12545 15860 15520
rect 16683 15560 16725 15569
rect 16683 15520 16684 15560
rect 16724 15520 16725 15560
rect 16683 15511 16725 15520
rect 16684 15426 16724 15511
rect 17644 15140 17684 17695
rect 17835 15728 17877 15737
rect 17835 15688 17836 15728
rect 17876 15688 17877 15728
rect 17835 15679 17877 15688
rect 17836 15594 17876 15679
rect 18124 15140 18164 23920
rect 19472 23456 19840 23465
rect 19512 23416 19554 23456
rect 19594 23416 19636 23456
rect 19676 23416 19718 23456
rect 19758 23416 19800 23456
rect 19472 23407 19840 23416
rect 21868 23129 21908 28792
rect 22059 28580 22101 28589
rect 22059 28540 22060 28580
rect 22100 28540 22101 28580
rect 22059 28531 22101 28540
rect 22060 28446 22100 28531
rect 22348 28328 22388 28337
rect 22348 27833 22388 28288
rect 22443 28328 22485 28337
rect 22443 28288 22444 28328
rect 22484 28288 22485 28328
rect 22443 28279 22485 28288
rect 22444 28194 22484 28279
rect 22540 28102 22580 28111
rect 22347 27824 22389 27833
rect 22347 27784 22348 27824
rect 22388 27784 22389 27824
rect 22347 27775 22389 27784
rect 22540 27749 22580 28062
rect 22539 27740 22581 27749
rect 22539 27700 22540 27740
rect 22580 27700 22581 27740
rect 22539 27691 22581 27700
rect 22636 26405 22676 31303
rect 23211 28328 23253 28337
rect 23211 28288 23212 28328
rect 23252 28288 23253 28328
rect 23211 28279 23253 28288
rect 23403 28328 23445 28337
rect 23403 28288 23404 28328
rect 23444 28288 23445 28328
rect 23403 28279 23445 28288
rect 23212 28244 23252 28279
rect 23212 28193 23252 28204
rect 23404 28085 23444 28279
rect 23500 28169 23540 35167
rect 33352 34796 33720 34805
rect 33392 34756 33434 34796
rect 33474 34756 33516 34796
rect 33556 34756 33598 34796
rect 33638 34756 33680 34796
rect 33352 34747 33720 34756
rect 48472 34796 48840 34805
rect 48512 34756 48554 34796
rect 48594 34756 48636 34796
rect 48676 34756 48718 34796
rect 48758 34756 48800 34796
rect 48472 34747 48840 34756
rect 63592 34796 63960 34805
rect 63632 34756 63674 34796
rect 63714 34756 63756 34796
rect 63796 34756 63838 34796
rect 63878 34756 63920 34796
rect 63592 34747 63960 34756
rect 78712 34796 79080 34805
rect 78752 34756 78794 34796
rect 78834 34756 78876 34796
rect 78916 34756 78958 34796
rect 78998 34756 79040 34796
rect 78712 34747 79080 34756
rect 93832 34796 94200 34805
rect 93872 34756 93914 34796
rect 93954 34756 93996 34796
rect 94036 34756 94078 34796
rect 94118 34756 94160 34796
rect 93832 34747 94200 34756
rect 29355 34376 29397 34385
rect 29355 34336 29356 34376
rect 29396 34336 29397 34376
rect 29355 34327 29397 34336
rect 29067 32864 29109 32873
rect 29067 32824 29068 32864
rect 29108 32824 29109 32864
rect 29067 32815 29109 32824
rect 27436 32192 27476 32201
rect 27051 31940 27093 31949
rect 27051 31900 27052 31940
rect 27092 31900 27093 31940
rect 27051 31891 27093 31900
rect 23787 31184 23829 31193
rect 23787 31144 23788 31184
rect 23828 31144 23829 31184
rect 23787 31135 23829 31144
rect 26764 31184 26804 31193
rect 23788 31050 23828 31135
rect 26764 30689 26804 31144
rect 26763 30680 26805 30689
rect 26763 30640 26764 30680
rect 26804 30640 26805 30680
rect 26763 30631 26805 30640
rect 23499 28160 23541 28169
rect 23499 28120 23500 28160
rect 23540 28120 23541 28160
rect 23499 28111 23541 28120
rect 26859 28160 26901 28169
rect 26859 28120 26860 28160
rect 26900 28120 26901 28160
rect 26859 28111 26901 28120
rect 23403 28076 23445 28085
rect 23403 28036 23404 28076
rect 23444 28036 23445 28076
rect 23403 28027 23445 28036
rect 23500 28026 23540 28111
rect 23307 27824 23349 27833
rect 26860 27824 26900 28111
rect 23307 27784 23308 27824
rect 23348 27784 23349 27824
rect 23307 27775 23349 27784
rect 26668 27784 26860 27824
rect 23308 27690 23348 27775
rect 23403 27740 23445 27749
rect 23403 27700 23404 27740
rect 23444 27700 23445 27740
rect 23403 27691 23445 27700
rect 26571 27740 26613 27749
rect 26571 27700 26572 27740
rect 26612 27700 26613 27740
rect 26571 27691 26613 27700
rect 23404 27656 23444 27691
rect 23404 27605 23444 27616
rect 26379 27656 26421 27665
rect 26379 27616 26380 27656
rect 26420 27616 26421 27656
rect 26379 27607 26421 27616
rect 23595 27404 23637 27413
rect 23595 27364 23596 27404
rect 23636 27364 23637 27404
rect 23595 27355 23637 27364
rect 23596 27270 23636 27355
rect 26380 26909 26420 27607
rect 26572 27606 26612 27691
rect 26668 27656 26708 27784
rect 26668 27607 26708 27616
rect 25803 26900 25845 26909
rect 25803 26860 25804 26900
rect 25844 26860 25845 26900
rect 25803 26851 25845 26860
rect 26379 26900 26421 26909
rect 26379 26860 26380 26900
rect 26420 26860 26421 26900
rect 26379 26851 26421 26860
rect 22635 26396 22677 26405
rect 22635 26356 22636 26396
rect 22676 26356 22677 26396
rect 22635 26347 22677 26356
rect 22636 24641 22676 26347
rect 25804 26312 25844 26851
rect 25804 26263 25844 26272
rect 26380 26144 26420 26153
rect 26380 26069 26420 26104
rect 26860 26069 26900 27784
rect 26955 27656 26997 27665
rect 26955 27616 26956 27656
rect 26996 27616 26997 27656
rect 26955 27607 26997 27616
rect 26956 27522 26996 27607
rect 25995 26060 26037 26069
rect 25995 26020 25996 26060
rect 26036 26020 26037 26060
rect 25995 26011 26037 26020
rect 26379 26060 26421 26069
rect 26379 26020 26380 26060
rect 26420 26020 26421 26060
rect 26379 26011 26421 26020
rect 26859 26060 26901 26069
rect 26859 26020 26860 26060
rect 26900 26020 26901 26060
rect 26859 26011 26901 26020
rect 25996 25926 26036 26011
rect 26380 25565 26420 26011
rect 26379 25556 26421 25565
rect 26379 25516 26380 25556
rect 26420 25516 26421 25556
rect 26379 25507 26421 25516
rect 22635 24632 22677 24641
rect 22635 24592 22636 24632
rect 22676 24592 22677 24632
rect 22635 24583 22677 24592
rect 23019 24632 23061 24641
rect 23019 24592 23020 24632
rect 23060 24592 23061 24632
rect 23019 24583 23061 24592
rect 23980 24632 24020 24641
rect 22636 24548 22676 24583
rect 22636 24498 22676 24508
rect 23020 24498 23060 24583
rect 19372 23120 19412 23129
rect 19180 23080 19372 23120
rect 18232 22700 18600 22709
rect 18272 22660 18314 22700
rect 18354 22660 18396 22700
rect 18436 22660 18478 22700
rect 18518 22660 18560 22700
rect 18232 22651 18600 22660
rect 18232 21188 18600 21197
rect 18272 21148 18314 21188
rect 18354 21148 18396 21188
rect 18436 21148 18478 21188
rect 18518 21148 18560 21188
rect 18232 21139 18600 21148
rect 19180 21020 19220 23080
rect 19372 23071 19412 23080
rect 19755 23120 19797 23129
rect 19755 23080 19756 23120
rect 19796 23080 19797 23120
rect 19755 23071 19797 23080
rect 20620 23120 20660 23129
rect 19756 22986 19796 23071
rect 19472 21944 19840 21953
rect 19512 21904 19554 21944
rect 19594 21904 19636 21944
rect 19676 21904 19718 21944
rect 19758 21904 19800 21944
rect 19472 21895 19840 21904
rect 19180 20971 19220 20980
rect 19276 20896 19508 20936
rect 18232 19676 18600 19685
rect 18272 19636 18314 19676
rect 18354 19636 18396 19676
rect 18436 19636 18478 19676
rect 18518 19636 18560 19676
rect 18232 19627 18600 19636
rect 19179 19340 19221 19349
rect 19179 19300 19180 19340
rect 19220 19300 19221 19340
rect 19179 19291 19221 19300
rect 19084 19256 19124 19267
rect 19084 19181 19124 19216
rect 19180 19206 19220 19291
rect 19083 19172 19125 19181
rect 19083 19132 19084 19172
rect 19124 19132 19125 19172
rect 19083 19123 19125 19132
rect 19276 19088 19316 20896
rect 19372 20768 19412 20777
rect 19372 19349 19412 20728
rect 19468 20768 19508 20896
rect 19468 20719 19508 20728
rect 19563 20768 19605 20777
rect 19563 20728 19564 20768
rect 19604 20728 19605 20768
rect 19563 20719 19605 20728
rect 20139 20768 20181 20777
rect 20139 20728 20140 20768
rect 20180 20728 20181 20768
rect 20139 20719 20181 20728
rect 19564 20634 19604 20719
rect 19472 20432 19840 20441
rect 19512 20392 19554 20432
rect 19594 20392 19636 20432
rect 19676 20392 19718 20432
rect 19758 20392 19800 20432
rect 19472 20383 19840 20392
rect 20140 20189 20180 20719
rect 20139 20180 20181 20189
rect 20139 20140 20140 20180
rect 20180 20140 20181 20180
rect 20139 20131 20181 20140
rect 19467 20096 19509 20105
rect 19467 20056 19468 20096
rect 19508 20056 19509 20096
rect 19467 20047 19509 20056
rect 19468 19517 19508 20047
rect 19467 19508 19509 19517
rect 19467 19468 19468 19508
rect 19508 19468 19509 19508
rect 19467 19459 19509 19468
rect 19371 19340 19413 19349
rect 19371 19300 19372 19340
rect 19412 19300 19413 19340
rect 19371 19291 19413 19300
rect 19468 19256 19508 19459
rect 19468 19207 19508 19216
rect 19659 19256 19701 19265
rect 19659 19216 19660 19256
rect 19700 19216 19701 19256
rect 19659 19207 19701 19216
rect 19660 19122 19700 19207
rect 19468 19088 19508 19097
rect 19276 19048 19468 19088
rect 18232 18164 18600 18173
rect 18272 18124 18314 18164
rect 18354 18124 18396 18164
rect 18436 18124 18478 18164
rect 18518 18124 18560 18164
rect 18232 18115 18600 18124
rect 19372 17753 19412 19048
rect 19468 19039 19508 19048
rect 19472 18920 19840 18929
rect 19512 18880 19554 18920
rect 19594 18880 19636 18920
rect 19676 18880 19718 18920
rect 19758 18880 19800 18920
rect 19472 18871 19840 18880
rect 19371 17744 19413 17753
rect 19371 17704 19372 17744
rect 19412 17704 19413 17744
rect 19371 17695 19413 17704
rect 19472 17408 19840 17417
rect 19512 17368 19554 17408
rect 19594 17368 19636 17408
rect 19676 17368 19718 17408
rect 19758 17368 19800 17408
rect 19472 17359 19840 17368
rect 18232 16652 18600 16661
rect 18272 16612 18314 16652
rect 18354 16612 18396 16652
rect 18436 16612 18478 16652
rect 18518 16612 18560 16652
rect 18232 16603 18600 16612
rect 19472 15896 19840 15905
rect 19512 15856 19554 15896
rect 19594 15856 19636 15896
rect 19676 15856 19718 15896
rect 19758 15856 19800 15896
rect 19472 15847 19840 15856
rect 18219 15728 18261 15737
rect 18219 15688 18220 15728
rect 18260 15688 18261 15728
rect 18219 15679 18261 15688
rect 18220 15594 18260 15679
rect 20620 15569 20660 23080
rect 21867 23120 21909 23129
rect 21867 23080 21868 23120
rect 21908 23080 21909 23120
rect 21867 23071 21909 23080
rect 21771 22868 21813 22877
rect 21771 22828 21772 22868
rect 21812 22828 21813 22868
rect 21771 22819 21813 22828
rect 21772 22734 21812 22819
rect 23403 22196 23445 22205
rect 23403 22156 23404 22196
rect 23444 22156 23445 22196
rect 23403 22147 23445 22156
rect 22635 20768 22677 20777
rect 22635 20728 22636 20768
rect 22676 20728 22677 20768
rect 22635 20719 22677 20728
rect 22732 20768 22772 20777
rect 22059 20348 22101 20357
rect 22059 20308 22060 20348
rect 22100 20308 22101 20348
rect 22059 20299 22101 20308
rect 22060 20264 22100 20299
rect 22060 20213 22100 20224
rect 21388 20105 21428 20190
rect 21771 20180 21813 20189
rect 21771 20140 21772 20180
rect 21812 20140 21813 20180
rect 21771 20131 21813 20140
rect 22347 20180 22389 20189
rect 22347 20140 22348 20180
rect 22388 20140 22389 20180
rect 22347 20131 22389 20140
rect 21100 20096 21140 20105
rect 21100 19349 21140 20056
rect 21196 20096 21236 20105
rect 21387 20096 21429 20105
rect 21236 20056 21332 20096
rect 21196 20047 21236 20056
rect 21099 19340 21141 19349
rect 21099 19300 21100 19340
rect 21140 19300 21141 19340
rect 21099 19291 21141 19300
rect 21100 18677 21140 19291
rect 21292 19265 21332 20056
rect 21387 20056 21388 20096
rect 21428 20056 21429 20096
rect 21387 20047 21429 20056
rect 21772 20096 21812 20131
rect 21772 20045 21812 20056
rect 21867 20096 21909 20105
rect 21867 20056 21868 20096
rect 21908 20056 21909 20096
rect 21867 20047 21909 20056
rect 21387 19928 21429 19937
rect 21387 19888 21388 19928
rect 21428 19888 21429 19928
rect 21387 19879 21429 19888
rect 21388 19794 21428 19879
rect 21291 19256 21333 19265
rect 21291 19216 21292 19256
rect 21332 19216 21333 19256
rect 21291 19207 21333 19216
rect 21099 18668 21141 18677
rect 21099 18628 21100 18668
rect 21140 18628 21141 18668
rect 21099 18619 21141 18628
rect 21292 17744 21332 19207
rect 21868 19172 21908 20047
rect 21772 19132 21908 19172
rect 21387 17996 21429 18005
rect 21387 17956 21388 17996
rect 21428 17956 21429 17996
rect 21387 17947 21429 17956
rect 21388 17862 21428 17947
rect 21292 17695 21332 17704
rect 21772 17744 21812 19132
rect 22252 18500 22292 18509
rect 21868 18124 22196 18164
rect 21868 17996 21908 18124
rect 21868 17947 21908 17956
rect 22059 17996 22101 18005
rect 22059 17956 22060 17996
rect 22100 17956 22101 17996
rect 22059 17947 22101 17956
rect 21772 17695 21812 17704
rect 22060 17072 22100 17947
rect 22060 17023 22100 17032
rect 22156 17744 22196 18124
rect 22252 18005 22292 18460
rect 22251 17996 22293 18005
rect 22251 17956 22252 17996
rect 22292 17956 22293 17996
rect 22251 17947 22293 17956
rect 18316 15560 18356 15569
rect 18316 15476 18356 15520
rect 18987 15560 19029 15569
rect 18987 15520 18988 15560
rect 19028 15520 19029 15560
rect 18987 15511 19029 15520
rect 20619 15560 20661 15569
rect 20619 15520 20620 15560
rect 20660 15520 20661 15560
rect 20619 15511 20661 15520
rect 18411 15476 18453 15485
rect 18316 15436 18412 15476
rect 18452 15436 18453 15476
rect 18411 15427 18453 15436
rect 18508 15401 18548 15486
rect 18892 15476 18932 15487
rect 18892 15401 18932 15436
rect 18507 15392 18549 15401
rect 18507 15352 18508 15392
rect 18548 15352 18549 15392
rect 18507 15343 18549 15352
rect 18891 15392 18933 15401
rect 18891 15352 18892 15392
rect 18932 15352 18933 15392
rect 18891 15343 18933 15352
rect 18699 15308 18741 15317
rect 18699 15268 18700 15308
rect 18740 15268 18741 15308
rect 18699 15259 18741 15268
rect 18700 15174 18740 15259
rect 17644 15100 17780 15140
rect 17740 12620 17780 15100
rect 17740 12571 17780 12580
rect 18028 15100 18164 15140
rect 18232 15140 18600 15149
rect 18892 15140 18932 15343
rect 18272 15100 18314 15140
rect 18354 15100 18396 15140
rect 18436 15100 18478 15140
rect 18518 15100 18560 15140
rect 15819 12536 15861 12545
rect 15819 12496 15820 12536
rect 15860 12496 15861 12536
rect 15819 12487 15861 12496
rect 3112 12116 3480 12125
rect 3152 12076 3194 12116
rect 3234 12076 3276 12116
rect 3316 12076 3358 12116
rect 3398 12076 3440 12116
rect 3112 12067 3480 12076
rect 4352 11360 4720 11369
rect 4392 11320 4434 11360
rect 4474 11320 4516 11360
rect 4556 11320 4598 11360
rect 4638 11320 4680 11360
rect 4352 11311 4720 11320
rect 18028 10949 18068 15100
rect 18232 15091 18600 15100
rect 18796 15100 18932 15140
rect 18232 13628 18600 13637
rect 18272 13588 18314 13628
rect 18354 13588 18396 13628
rect 18436 13588 18478 13628
rect 18518 13588 18560 13628
rect 18232 13579 18600 13588
rect 18123 12536 18165 12545
rect 18123 12496 18124 12536
rect 18164 12496 18165 12536
rect 18123 12487 18165 12496
rect 18124 12402 18164 12487
rect 18232 12116 18600 12125
rect 18272 12076 18314 12116
rect 18354 12076 18396 12116
rect 18436 12076 18478 12116
rect 18518 12076 18560 12116
rect 18232 12067 18600 12076
rect 18027 10940 18069 10949
rect 18027 10900 18028 10940
rect 18068 10900 18069 10940
rect 18027 10891 18069 10900
rect 3112 10604 3480 10613
rect 3152 10564 3194 10604
rect 3234 10564 3276 10604
rect 3316 10564 3358 10604
rect 3398 10564 3440 10604
rect 3112 10555 3480 10564
rect 18232 10604 18600 10613
rect 18272 10564 18314 10604
rect 18354 10564 18396 10604
rect 18436 10564 18478 10604
rect 18518 10564 18560 10604
rect 18232 10555 18600 10564
rect 4352 9848 4720 9857
rect 4392 9808 4434 9848
rect 4474 9808 4516 9848
rect 4556 9808 4598 9848
rect 4638 9808 4680 9848
rect 4352 9799 4720 9808
rect 3112 9092 3480 9101
rect 3152 9052 3194 9092
rect 3234 9052 3276 9092
rect 3316 9052 3358 9092
rect 3398 9052 3440 9092
rect 3112 9043 3480 9052
rect 18232 9092 18600 9101
rect 18272 9052 18314 9092
rect 18354 9052 18396 9092
rect 18436 9052 18478 9092
rect 18518 9052 18560 9092
rect 18232 9043 18600 9052
rect 4352 8336 4720 8345
rect 4392 8296 4434 8336
rect 4474 8296 4516 8336
rect 4556 8296 4598 8336
rect 4638 8296 4680 8336
rect 4352 8287 4720 8296
rect 3112 7580 3480 7589
rect 3152 7540 3194 7580
rect 3234 7540 3276 7580
rect 3316 7540 3358 7580
rect 3398 7540 3440 7580
rect 3112 7531 3480 7540
rect 18232 7580 18600 7589
rect 18272 7540 18314 7580
rect 18354 7540 18396 7580
rect 18436 7540 18478 7580
rect 18518 7540 18560 7580
rect 18232 7531 18600 7540
rect 4352 6824 4720 6833
rect 4392 6784 4434 6824
rect 4474 6784 4516 6824
rect 4556 6784 4598 6824
rect 4638 6784 4680 6824
rect 4352 6775 4720 6784
rect 18796 6320 18836 15100
rect 18988 12536 19028 15511
rect 22156 15140 22196 17704
rect 22348 17744 22388 20131
rect 22539 19172 22581 19181
rect 22539 19132 22540 19172
rect 22580 19132 22581 19172
rect 22539 19123 22581 19132
rect 22443 18668 22485 18677
rect 22443 18628 22444 18668
rect 22484 18628 22485 18668
rect 22443 18619 22485 18628
rect 22444 18584 22484 18619
rect 22444 18533 22484 18544
rect 22443 18332 22485 18341
rect 22443 18292 22444 18332
rect 22484 18292 22485 18332
rect 22443 18283 22485 18292
rect 22444 18198 22484 18283
rect 22348 17695 22388 17704
rect 22540 17744 22580 19123
rect 22636 18341 22676 20719
rect 22732 20357 22772 20728
rect 22828 20768 22868 20777
rect 22731 20348 22773 20357
rect 22731 20308 22732 20348
rect 22772 20308 22773 20348
rect 22731 20299 22773 20308
rect 22828 20180 22868 20728
rect 23116 20768 23156 20777
rect 22923 20684 22965 20693
rect 22923 20644 22924 20684
rect 22964 20644 22965 20684
rect 22923 20635 22965 20644
rect 22924 20550 22964 20635
rect 23116 20273 23156 20728
rect 23211 20768 23253 20777
rect 23211 20728 23212 20768
rect 23252 20728 23253 20768
rect 23211 20719 23253 20728
rect 23308 20768 23348 20777
rect 23212 20634 23252 20719
rect 23115 20264 23157 20273
rect 23115 20224 23116 20264
rect 23156 20224 23157 20264
rect 23115 20215 23157 20224
rect 22732 20140 22868 20180
rect 22732 19937 22772 20140
rect 23212 20096 23252 20105
rect 22828 20056 23212 20096
rect 22828 20012 22868 20056
rect 23212 20047 23252 20056
rect 22828 19963 22868 19972
rect 23308 19937 23348 20728
rect 23404 20768 23444 22147
rect 23980 21533 24020 24592
rect 25419 23876 25461 23885
rect 25419 23836 25420 23876
rect 25460 23836 25461 23876
rect 25419 23827 25461 23836
rect 24555 23120 24597 23129
rect 24555 23080 24556 23120
rect 24596 23080 24597 23120
rect 24555 23071 24597 23080
rect 24556 22280 24596 23071
rect 24556 22231 24596 22240
rect 25420 22280 25460 23827
rect 26571 22364 26613 22373
rect 26571 22324 26572 22364
rect 26612 22324 26613 22364
rect 26571 22315 26613 22324
rect 25420 22231 25460 22240
rect 26572 22230 26612 22315
rect 24171 22196 24213 22205
rect 24171 22156 24172 22196
rect 24212 22156 24213 22196
rect 24171 22147 24213 22156
rect 24172 22062 24212 22147
rect 23979 21524 24021 21533
rect 23979 21484 23980 21524
rect 24020 21484 24021 21524
rect 23979 21475 24021 21484
rect 24171 21524 24213 21533
rect 24171 21484 24172 21524
rect 24212 21484 24213 21524
rect 24171 21475 24213 21484
rect 23404 20719 23444 20728
rect 23499 20180 23541 20189
rect 23499 20140 23500 20180
rect 23540 20140 23541 20180
rect 23499 20131 23541 20140
rect 22731 19928 22773 19937
rect 22731 19888 22732 19928
rect 22772 19888 22773 19928
rect 22731 19879 22773 19888
rect 23307 19928 23349 19937
rect 23307 19888 23308 19928
rect 23348 19888 23349 19928
rect 23307 19879 23349 19888
rect 23500 19265 23540 20131
rect 24172 20096 24212 21475
rect 24172 20047 24212 20056
rect 23692 19844 23732 19853
rect 23732 19804 23828 19844
rect 23692 19795 23732 19804
rect 23499 19256 23541 19265
rect 23499 19216 23500 19256
rect 23540 19216 23541 19256
rect 23499 19207 23541 19216
rect 22731 18500 22773 18509
rect 22731 18460 22732 18500
rect 22772 18460 22773 18500
rect 22731 18451 22773 18460
rect 22635 18332 22677 18341
rect 22635 18292 22636 18332
rect 22676 18292 22677 18332
rect 22635 18283 22677 18292
rect 22732 17753 22772 18451
rect 22828 17912 22868 17921
rect 22868 17872 22964 17912
rect 22828 17863 22868 17872
rect 22251 17660 22293 17669
rect 22251 17620 22252 17660
rect 22292 17620 22293 17660
rect 22251 17611 22293 17620
rect 22252 17492 22292 17611
rect 22252 17452 22388 17492
rect 22251 17072 22293 17081
rect 22251 17032 22252 17072
rect 22292 17032 22293 17072
rect 22251 17023 22293 17032
rect 22348 17072 22388 17452
rect 22540 17081 22580 17704
rect 22731 17744 22773 17753
rect 22731 17704 22732 17744
rect 22772 17704 22773 17744
rect 22731 17695 22773 17704
rect 22828 17744 22868 17755
rect 22924 17753 22964 17872
rect 22732 17610 22772 17695
rect 22828 17669 22868 17704
rect 22923 17744 22965 17753
rect 22923 17704 22924 17744
rect 22964 17704 22965 17744
rect 22923 17695 22965 17704
rect 22827 17660 22869 17669
rect 22827 17620 22828 17660
rect 22868 17620 22869 17660
rect 22827 17611 22869 17620
rect 22348 17023 22388 17032
rect 22539 17072 22581 17081
rect 22539 17032 22540 17072
rect 22580 17032 22581 17072
rect 22539 17023 22581 17032
rect 22252 16938 22292 17023
rect 23019 16988 23061 16997
rect 23019 16948 23020 16988
rect 23060 16948 23061 16988
rect 23019 16939 23061 16948
rect 22348 16904 22388 16913
rect 22388 16864 22676 16904
rect 22348 16855 22388 16864
rect 22156 15100 22580 15140
rect 19472 14384 19840 14393
rect 19512 14344 19554 14384
rect 19594 14344 19636 14384
rect 19676 14344 19718 14384
rect 19758 14344 19800 14384
rect 19472 14335 19840 14344
rect 19472 12872 19840 12881
rect 19512 12832 19554 12872
rect 19594 12832 19636 12872
rect 19676 12832 19718 12872
rect 19758 12832 19800 12872
rect 19472 12823 19840 12832
rect 18988 12487 19028 12496
rect 20139 12284 20181 12293
rect 20139 12244 20140 12284
rect 20180 12244 20181 12284
rect 20139 12235 20181 12244
rect 20140 12150 20180 12235
rect 22540 11696 22580 15100
rect 22636 14720 22676 16864
rect 22636 14671 22676 14680
rect 23020 14720 23060 16939
rect 23788 15569 23828 19804
rect 26475 18752 26517 18761
rect 26475 18712 26476 18752
rect 26516 18712 26517 18752
rect 26475 18703 26517 18712
rect 26091 18668 26133 18677
rect 26091 18628 26092 18668
rect 26132 18628 26133 18668
rect 26091 18619 26133 18628
rect 26092 18584 26132 18619
rect 26092 18533 26132 18544
rect 26476 18584 26516 18703
rect 26187 18500 26229 18509
rect 26187 18460 26188 18500
rect 26228 18460 26229 18500
rect 26187 18451 26229 18460
rect 26379 18500 26421 18509
rect 26379 18460 26380 18500
rect 26420 18460 26421 18500
rect 26379 18451 26421 18460
rect 26188 18366 26228 18451
rect 26284 18416 26324 18425
rect 26284 17753 26324 18376
rect 26380 18366 26420 18451
rect 26476 18341 26516 18544
rect 26475 18332 26517 18341
rect 26475 18292 26476 18332
rect 26516 18292 26517 18332
rect 26475 18283 26517 18292
rect 26283 17744 26325 17753
rect 26283 17704 26284 17744
rect 26324 17704 26325 17744
rect 26283 17695 26325 17704
rect 26763 17744 26805 17753
rect 26763 17704 26764 17744
rect 26804 17704 26805 17744
rect 26763 17695 26805 17704
rect 26764 17610 26804 17695
rect 23787 15560 23829 15569
rect 23787 15520 23788 15560
rect 23828 15520 23829 15560
rect 23787 15511 23829 15520
rect 25035 15560 25077 15569
rect 25035 15520 25036 15560
rect 25076 15520 25077 15560
rect 25035 15511 25077 15520
rect 23020 12545 23060 14680
rect 23788 14720 23828 15511
rect 25036 14972 25076 15511
rect 25036 14923 25076 14932
rect 23884 14720 23924 14729
rect 23788 14680 23884 14720
rect 23019 12536 23061 12545
rect 23019 12496 23020 12536
rect 23060 12496 23061 12536
rect 23019 12487 23061 12496
rect 22540 11647 22580 11656
rect 22924 11696 22964 11705
rect 23020 11696 23060 12487
rect 22964 11656 23060 11696
rect 23788 11696 23828 14680
rect 23884 14671 23924 14680
rect 26955 13208 26997 13217
rect 26955 13168 26956 13208
rect 26996 13168 26997 13208
rect 26955 13159 26997 13168
rect 26859 12788 26901 12797
rect 26859 12748 26860 12788
rect 26900 12748 26901 12788
rect 26859 12739 26901 12748
rect 26571 12704 26613 12713
rect 26571 12664 26572 12704
rect 26612 12664 26613 12704
rect 26571 12655 26613 12664
rect 26475 12620 26517 12629
rect 26475 12580 26476 12620
rect 26516 12580 26517 12620
rect 26475 12571 26517 12580
rect 26380 12536 26420 12545
rect 26380 11957 26420 12496
rect 26476 12486 26516 12571
rect 26572 12536 26612 12655
rect 26860 12620 26900 12739
rect 26956 12713 26996 13159
rect 26955 12704 26997 12713
rect 26955 12664 26956 12704
rect 26996 12664 26997 12704
rect 26955 12655 26997 12664
rect 26860 12571 26900 12580
rect 26572 12487 26612 12496
rect 26764 12536 26804 12545
rect 26764 12293 26804 12496
rect 26956 12536 26996 12655
rect 26956 12487 26996 12496
rect 26763 12284 26805 12293
rect 26763 12244 26764 12284
rect 26804 12244 26805 12284
rect 26763 12235 26805 12244
rect 24939 11948 24981 11957
rect 24939 11908 24940 11948
rect 24980 11908 24981 11948
rect 24939 11899 24981 11908
rect 26379 11948 26421 11957
rect 26379 11908 26380 11948
rect 26420 11908 26421 11948
rect 26379 11899 26421 11908
rect 24940 11814 24980 11899
rect 22924 11647 22964 11656
rect 23788 11647 23828 11656
rect 19472 11360 19840 11369
rect 19512 11320 19554 11360
rect 19594 11320 19636 11360
rect 19676 11320 19718 11360
rect 19758 11320 19800 11360
rect 19472 11311 19840 11320
rect 19472 9848 19840 9857
rect 19512 9808 19554 9848
rect 19594 9808 19636 9848
rect 19676 9808 19718 9848
rect 19758 9808 19800 9848
rect 19472 9799 19840 9808
rect 27052 9437 27092 31891
rect 27339 31184 27381 31193
rect 27339 31144 27340 31184
rect 27380 31144 27381 31184
rect 27339 31135 27381 31144
rect 27244 30680 27284 30689
rect 27147 28328 27189 28337
rect 27147 28288 27148 28328
rect 27188 28288 27189 28328
rect 27147 28279 27189 28288
rect 27148 27740 27188 28279
rect 27148 27691 27188 27700
rect 27244 26144 27284 30640
rect 27340 30596 27380 31135
rect 27340 30547 27380 30556
rect 27436 30512 27476 32152
rect 27531 31940 27573 31949
rect 27531 31900 27532 31940
rect 27572 31900 27573 31940
rect 27531 31891 27573 31900
rect 27532 31806 27572 31891
rect 27915 31352 27957 31361
rect 27915 31312 27916 31352
rect 27956 31312 27957 31352
rect 27915 31303 27957 31312
rect 28780 31352 28820 31363
rect 27916 31218 27956 31303
rect 28780 31277 28820 31312
rect 28779 31268 28821 31277
rect 28779 31228 28780 31268
rect 28820 31228 28821 31268
rect 28779 31219 28821 31228
rect 27627 30680 27669 30689
rect 27627 30640 27628 30680
rect 27668 30640 27669 30680
rect 27627 30631 27669 30640
rect 27436 30463 27476 30472
rect 27532 30596 27572 30605
rect 27532 28421 27572 30556
rect 27628 30546 27668 30631
rect 28780 30605 28820 31219
rect 28779 30596 28821 30605
rect 28779 30556 28780 30596
rect 28820 30556 28821 30596
rect 28779 30547 28821 30556
rect 28299 30260 28341 30269
rect 28299 30220 28300 30260
rect 28340 30220 28341 30260
rect 28299 30211 28341 30220
rect 28203 28496 28245 28505
rect 28203 28456 28204 28496
rect 28244 28456 28245 28496
rect 28203 28447 28245 28456
rect 28300 28496 28340 30211
rect 29068 28832 29108 32815
rect 29164 31268 29204 31277
rect 29164 30269 29204 31228
rect 29163 30260 29205 30269
rect 29163 30220 29164 30260
rect 29204 30220 29205 30260
rect 29163 30211 29205 30220
rect 29068 28792 29204 28832
rect 28300 28447 28340 28456
rect 28779 28496 28821 28505
rect 28779 28456 28780 28496
rect 28820 28456 28821 28496
rect 28779 28447 28821 28456
rect 27531 28412 27573 28421
rect 27531 28372 27532 28412
rect 27572 28372 27573 28412
rect 27531 28363 27573 28372
rect 28204 28412 28244 28447
rect 27244 22541 27284 26104
rect 27532 24557 27572 28363
rect 28204 28361 28244 28372
rect 28396 28412 28436 28421
rect 28107 28328 28149 28337
rect 28107 28288 28108 28328
rect 28148 28288 28149 28328
rect 28107 28279 28149 28288
rect 28011 28244 28053 28253
rect 28011 28204 28012 28244
rect 28052 28204 28053 28244
rect 28011 28195 28053 28204
rect 28012 25145 28052 28195
rect 28108 28194 28148 28279
rect 28299 27824 28341 27833
rect 28299 27784 28300 27824
rect 28340 27784 28341 27824
rect 28299 27775 28341 27784
rect 28107 27488 28149 27497
rect 28107 27448 28108 27488
rect 28148 27448 28149 27488
rect 28107 27439 28149 27448
rect 28108 25976 28148 27439
rect 28300 26312 28340 27775
rect 28396 27749 28436 28372
rect 28780 28362 28820 28447
rect 28492 28328 28532 28337
rect 28492 28169 28532 28288
rect 29068 28328 29108 28337
rect 28491 28160 28533 28169
rect 28491 28120 28492 28160
rect 28532 28120 28533 28160
rect 28491 28111 28533 28120
rect 28395 27740 28437 27749
rect 28395 27700 28396 27740
rect 28436 27700 28437 27740
rect 28395 27691 28437 27700
rect 29068 27152 29108 28288
rect 29164 28328 29204 28792
rect 29164 27581 29204 28288
rect 29356 28328 29396 34327
rect 34592 34040 34960 34049
rect 34632 34000 34674 34040
rect 34714 34000 34756 34040
rect 34796 34000 34838 34040
rect 34878 34000 34920 34040
rect 34592 33991 34960 34000
rect 49712 34040 50080 34049
rect 49752 34000 49794 34040
rect 49834 34000 49876 34040
rect 49916 34000 49958 34040
rect 49998 34000 50040 34040
rect 49712 33991 50080 34000
rect 64832 34040 65200 34049
rect 64872 34000 64914 34040
rect 64954 34000 64996 34040
rect 65036 34000 65078 34040
rect 65118 34000 65160 34040
rect 64832 33991 65200 34000
rect 79952 34040 80320 34049
rect 79992 34000 80034 34040
rect 80074 34000 80116 34040
rect 80156 34000 80198 34040
rect 80238 34000 80280 34040
rect 79952 33991 80320 34000
rect 95072 34040 95440 34049
rect 95112 34000 95154 34040
rect 95194 34000 95236 34040
rect 95276 34000 95318 34040
rect 95358 34000 95400 34040
rect 95072 33991 95440 34000
rect 29643 33704 29685 33713
rect 29643 33664 29644 33704
rect 29684 33664 29685 33704
rect 29643 33655 29685 33664
rect 29452 28328 29492 28337
rect 29644 28328 29684 33655
rect 33352 33284 33720 33293
rect 33392 33244 33434 33284
rect 33474 33244 33516 33284
rect 33556 33244 33598 33284
rect 33638 33244 33680 33284
rect 33352 33235 33720 33244
rect 48472 33284 48840 33293
rect 48512 33244 48554 33284
rect 48594 33244 48636 33284
rect 48676 33244 48718 33284
rect 48758 33244 48800 33284
rect 48472 33235 48840 33244
rect 63592 33284 63960 33293
rect 63632 33244 63674 33284
rect 63714 33244 63756 33284
rect 63796 33244 63838 33284
rect 63878 33244 63920 33284
rect 63592 33235 63960 33244
rect 78712 33284 79080 33293
rect 78752 33244 78794 33284
rect 78834 33244 78876 33284
rect 78916 33244 78958 33284
rect 78998 33244 79040 33284
rect 78712 33235 79080 33244
rect 93832 33284 94200 33293
rect 93872 33244 93914 33284
rect 93954 33244 93996 33284
rect 94036 33244 94078 33284
rect 94118 33244 94160 33284
rect 93832 33235 94200 33244
rect 34592 32528 34960 32537
rect 34632 32488 34674 32528
rect 34714 32488 34756 32528
rect 34796 32488 34838 32528
rect 34878 32488 34920 32528
rect 34592 32479 34960 32488
rect 49712 32528 50080 32537
rect 49752 32488 49794 32528
rect 49834 32488 49876 32528
rect 49916 32488 49958 32528
rect 49998 32488 50040 32528
rect 49712 32479 50080 32488
rect 64832 32528 65200 32537
rect 64872 32488 64914 32528
rect 64954 32488 64996 32528
rect 65036 32488 65078 32528
rect 65118 32488 65160 32528
rect 64832 32479 65200 32488
rect 79952 32528 80320 32537
rect 79992 32488 80034 32528
rect 80074 32488 80116 32528
rect 80156 32488 80198 32528
rect 80238 32488 80280 32528
rect 79952 32479 80320 32488
rect 95072 32528 95440 32537
rect 95112 32488 95154 32528
rect 95194 32488 95236 32528
rect 95276 32488 95318 32528
rect 95358 32488 95400 32528
rect 95072 32479 95440 32488
rect 33352 31772 33720 31781
rect 33392 31732 33434 31772
rect 33474 31732 33516 31772
rect 33556 31732 33598 31772
rect 33638 31732 33680 31772
rect 33352 31723 33720 31732
rect 48472 31772 48840 31781
rect 48512 31732 48554 31772
rect 48594 31732 48636 31772
rect 48676 31732 48718 31772
rect 48758 31732 48800 31772
rect 48472 31723 48840 31732
rect 63592 31772 63960 31781
rect 63632 31732 63674 31772
rect 63714 31732 63756 31772
rect 63796 31732 63838 31772
rect 63878 31732 63920 31772
rect 63592 31723 63960 31732
rect 78712 31772 79080 31781
rect 78752 31732 78794 31772
rect 78834 31732 78876 31772
rect 78916 31732 78958 31772
rect 78998 31732 79040 31772
rect 78712 31723 79080 31732
rect 93832 31772 94200 31781
rect 93872 31732 93914 31772
rect 93954 31732 93996 31772
rect 94036 31732 94078 31772
rect 94118 31732 94160 31772
rect 93832 31723 94200 31732
rect 34592 31016 34960 31025
rect 34632 30976 34674 31016
rect 34714 30976 34756 31016
rect 34796 30976 34838 31016
rect 34878 30976 34920 31016
rect 34592 30967 34960 30976
rect 49712 31016 50080 31025
rect 49752 30976 49794 31016
rect 49834 30976 49876 31016
rect 49916 30976 49958 31016
rect 49998 30976 50040 31016
rect 49712 30967 50080 30976
rect 64832 31016 65200 31025
rect 64872 30976 64914 31016
rect 64954 30976 64996 31016
rect 65036 30976 65078 31016
rect 65118 30976 65160 31016
rect 64832 30967 65200 30976
rect 79952 31016 80320 31025
rect 79992 30976 80034 31016
rect 80074 30976 80116 31016
rect 80156 30976 80198 31016
rect 80238 30976 80280 31016
rect 79952 30967 80320 30976
rect 95072 31016 95440 31025
rect 95112 30976 95154 31016
rect 95194 30976 95236 31016
rect 95276 30976 95318 31016
rect 95358 30976 95400 31016
rect 95072 30967 95440 30976
rect 32716 30680 32756 30689
rect 32716 30269 32756 30640
rect 32811 30680 32853 30689
rect 32811 30640 32812 30680
rect 32852 30640 32853 30680
rect 32811 30631 32853 30640
rect 33100 30680 33140 30691
rect 31275 30260 31317 30269
rect 31275 30220 31276 30260
rect 31316 30220 31317 30260
rect 31275 30211 31317 30220
rect 32715 30260 32757 30269
rect 32715 30220 32716 30260
rect 32756 30220 32757 30260
rect 32715 30211 32757 30220
rect 31276 29336 31316 30211
rect 31276 29287 31316 29296
rect 31180 29168 31220 29177
rect 31180 28337 31220 29128
rect 29356 28288 29452 28328
rect 29260 28102 29300 28111
rect 29260 27656 29300 28062
rect 29356 27740 29396 28288
rect 29452 28279 29492 28288
rect 29548 28288 29644 28328
rect 29451 28160 29493 28169
rect 29451 28120 29452 28160
rect 29492 28120 29493 28160
rect 29451 28111 29493 28120
rect 29452 28026 29492 28111
rect 29451 27740 29493 27749
rect 29356 27700 29452 27740
rect 29492 27700 29493 27740
rect 29451 27691 29493 27700
rect 29548 27656 29588 28288
rect 29644 28279 29684 28288
rect 29740 28328 29780 28337
rect 31179 28328 31221 28337
rect 29780 28288 29972 28328
rect 29740 28279 29780 28288
rect 29260 27616 29396 27656
rect 29163 27572 29205 27581
rect 29163 27532 29164 27572
rect 29204 27532 29205 27572
rect 29163 27523 29205 27532
rect 29259 27488 29301 27497
rect 29259 27448 29260 27488
rect 29300 27448 29301 27488
rect 29259 27439 29301 27448
rect 29356 27446 29396 27616
rect 29451 27572 29493 27581
rect 29451 27532 29452 27572
rect 29492 27532 29493 27572
rect 29451 27523 29493 27532
rect 29260 27354 29300 27439
rect 29355 27406 29356 27413
rect 29452 27438 29492 27523
rect 29396 27406 29397 27413
rect 29355 27404 29397 27406
rect 29355 27364 29356 27404
rect 29396 27364 29397 27404
rect 29355 27355 29397 27364
rect 29356 27311 29396 27355
rect 29068 27112 29492 27152
rect 29452 27068 29492 27112
rect 29452 27019 29492 27028
rect 29548 26984 29588 27616
rect 29643 27656 29685 27665
rect 29643 27607 29644 27656
rect 29684 27607 29685 27656
rect 29644 27152 29684 27600
rect 29644 27112 29780 27152
rect 29644 26984 29684 26993
rect 29548 26944 29644 26984
rect 29644 26935 29684 26944
rect 29644 26816 29684 26825
rect 29740 26816 29780 27112
rect 29932 27068 29972 28288
rect 31179 28288 31180 28328
rect 31220 28288 31221 28328
rect 31179 28279 31221 28288
rect 30027 27572 30069 27581
rect 30027 27532 30028 27572
rect 30068 27532 30069 27572
rect 30027 27523 30069 27532
rect 29932 27019 29972 27028
rect 29684 26776 29780 26816
rect 30028 26816 30068 27523
rect 30123 27404 30165 27413
rect 30123 27364 30124 27404
rect 30164 27364 30165 27404
rect 30123 27355 30165 27364
rect 30124 26984 30164 27355
rect 30164 26944 30260 26984
rect 30124 26935 30164 26944
rect 30124 26816 30164 26825
rect 30028 26776 30124 26816
rect 29644 26767 29684 26776
rect 30124 26767 30164 26776
rect 28300 26263 28340 26272
rect 28300 26144 28340 26153
rect 28203 26060 28245 26069
rect 28203 26020 28204 26060
rect 28244 26020 28245 26060
rect 28203 26011 28245 26020
rect 28108 25927 28148 25936
rect 28204 25926 28244 26011
rect 28203 25556 28245 25565
rect 28203 25516 28204 25556
rect 28244 25516 28245 25556
rect 28203 25507 28245 25516
rect 28204 25422 28244 25507
rect 28300 25304 28340 26104
rect 28396 26144 28436 26153
rect 28436 26104 28628 26144
rect 28396 26095 28436 26104
rect 28395 25304 28437 25313
rect 28300 25264 28396 25304
rect 28436 25264 28437 25304
rect 28395 25255 28437 25264
rect 28396 25170 28436 25255
rect 28011 25136 28053 25145
rect 28011 25096 28012 25136
rect 28052 25096 28053 25136
rect 28011 25087 28053 25096
rect 28491 25136 28533 25145
rect 28491 25096 28492 25136
rect 28532 25096 28533 25136
rect 28491 25087 28533 25096
rect 27531 24548 27573 24557
rect 27531 24508 27532 24548
rect 27572 24508 27573 24548
rect 27531 24499 27573 24508
rect 28492 23717 28532 25087
rect 28588 23960 28628 26104
rect 29259 25304 29301 25313
rect 29259 25264 29260 25304
rect 29300 25264 29301 25304
rect 29259 25255 29301 25264
rect 30027 25304 30069 25313
rect 30027 25264 30028 25304
rect 30068 25264 30069 25304
rect 30027 25255 30069 25264
rect 28876 23960 28916 23969
rect 28588 23920 28876 23960
rect 28491 23708 28533 23717
rect 28491 23668 28492 23708
rect 28532 23668 28533 23708
rect 28491 23659 28533 23668
rect 28588 23288 28628 23920
rect 28492 23248 28628 23288
rect 27243 22532 27285 22541
rect 27243 22492 27244 22532
rect 27284 22492 27285 22532
rect 27243 22483 27285 22492
rect 28492 22280 28532 23248
rect 28588 23120 28628 23129
rect 28588 22877 28628 23080
rect 28684 23120 28724 23129
rect 28587 22868 28629 22877
rect 28587 22828 28588 22868
rect 28628 22828 28629 22868
rect 28587 22819 28629 22828
rect 28684 22457 28724 23080
rect 28876 23120 28916 23920
rect 28972 23792 29012 23801
rect 28972 23717 29012 23752
rect 28971 23708 29013 23717
rect 28971 23668 28972 23708
rect 29012 23668 29013 23708
rect 28971 23659 29013 23668
rect 28972 23288 29012 23659
rect 28972 23248 29108 23288
rect 28876 23071 28916 23080
rect 28876 22868 28916 22877
rect 28876 22625 28916 22828
rect 28875 22616 28917 22625
rect 28875 22576 28876 22616
rect 28916 22576 28917 22616
rect 28875 22567 28917 22576
rect 28683 22448 28725 22457
rect 28683 22408 28684 22448
rect 28724 22408 28725 22448
rect 28683 22399 28725 22408
rect 28875 22448 28917 22457
rect 28875 22408 28876 22448
rect 28916 22408 28917 22448
rect 28875 22399 28917 22408
rect 28779 22364 28821 22373
rect 28779 22324 28780 22364
rect 28820 22324 28821 22364
rect 28779 22315 28821 22324
rect 28684 22280 28724 22289
rect 28492 22240 28684 22280
rect 28684 22231 28724 22240
rect 28780 22280 28820 22315
rect 28780 22229 28820 22240
rect 28876 22280 28916 22399
rect 28876 22231 28916 22240
rect 28972 22112 29012 22121
rect 28876 22072 28972 22112
rect 28395 21608 28437 21617
rect 28395 21568 28396 21608
rect 28436 21568 28437 21608
rect 28395 21559 28437 21568
rect 28396 21474 28436 21559
rect 28876 20861 28916 22072
rect 28972 22063 29012 22072
rect 29068 20936 29108 23248
rect 29163 22448 29205 22457
rect 29163 22408 29164 22448
rect 29204 22408 29205 22448
rect 29163 22399 29205 22408
rect 29164 22314 29204 22399
rect 29260 22280 29300 25255
rect 29644 24800 29684 24809
rect 29644 23717 29684 24760
rect 29836 24716 29876 24725
rect 29836 24557 29876 24676
rect 30028 24632 30068 25255
rect 30028 24583 30068 24592
rect 29835 24548 29877 24557
rect 29835 24508 29836 24548
rect 29876 24508 29877 24548
rect 29835 24499 29877 24508
rect 30220 23960 30260 26944
rect 30124 23920 30260 23960
rect 30124 23801 30164 23920
rect 32812 23885 32852 30631
rect 33100 30605 33140 30640
rect 33963 30680 34005 30689
rect 33963 30640 33964 30680
rect 34004 30640 34005 30680
rect 33963 30631 34005 30640
rect 33099 30596 33141 30605
rect 33099 30556 33100 30596
rect 33140 30556 33141 30596
rect 33099 30547 33141 30556
rect 33964 30546 34004 30631
rect 34347 30596 34389 30605
rect 34347 30556 34348 30596
rect 34388 30556 34389 30596
rect 34347 30547 34389 30556
rect 33352 30260 33720 30269
rect 33392 30220 33434 30260
rect 33474 30220 33516 30260
rect 33556 30220 33598 30260
rect 33638 30220 33680 30260
rect 33352 30211 33720 30220
rect 33352 28748 33720 28757
rect 33392 28708 33434 28748
rect 33474 28708 33516 28748
rect 33556 28708 33598 28748
rect 33638 28708 33680 28748
rect 33352 28699 33720 28708
rect 33352 27236 33720 27245
rect 33392 27196 33434 27236
rect 33474 27196 33516 27236
rect 33556 27196 33598 27236
rect 33638 27196 33680 27236
rect 33352 27187 33720 27196
rect 34348 26144 34388 30547
rect 35115 30428 35157 30437
rect 35115 30388 35116 30428
rect 35156 30388 35157 30428
rect 35115 30379 35157 30388
rect 35595 30428 35637 30437
rect 35595 30388 35596 30428
rect 35636 30388 35637 30428
rect 35595 30379 35637 30388
rect 35116 30294 35156 30379
rect 34592 29504 34960 29513
rect 34632 29464 34674 29504
rect 34714 29464 34756 29504
rect 34796 29464 34838 29504
rect 34878 29464 34920 29504
rect 34592 29455 34960 29464
rect 35596 29168 35636 30379
rect 48472 30260 48840 30269
rect 48512 30220 48554 30260
rect 48594 30220 48636 30260
rect 48676 30220 48718 30260
rect 48758 30220 48800 30260
rect 48472 30211 48840 30220
rect 63592 30260 63960 30269
rect 63632 30220 63674 30260
rect 63714 30220 63756 30260
rect 63796 30220 63838 30260
rect 63878 30220 63920 30260
rect 63592 30211 63960 30220
rect 78712 30260 79080 30269
rect 78752 30220 78794 30260
rect 78834 30220 78876 30260
rect 78916 30220 78958 30260
rect 78998 30220 79040 30260
rect 78712 30211 79080 30220
rect 93832 30260 94200 30269
rect 93872 30220 93914 30260
rect 93954 30220 93996 30260
rect 94036 30220 94078 30260
rect 94118 30220 94160 30260
rect 93832 30211 94200 30220
rect 36460 29840 36500 29849
rect 35596 29119 35636 29128
rect 35980 29168 36020 29177
rect 36020 29128 36116 29168
rect 35980 29119 36020 29128
rect 35692 29084 35732 29093
rect 34592 27992 34960 28001
rect 34632 27952 34674 27992
rect 34714 27952 34756 27992
rect 34796 27952 34838 27992
rect 34878 27952 34920 27992
rect 34592 27943 34960 27952
rect 34923 27320 34965 27329
rect 34923 27280 34924 27320
rect 34964 27280 34965 27320
rect 34923 27271 34965 27280
rect 34924 26816 34964 27271
rect 35692 26900 35732 29044
rect 35884 29084 35924 29093
rect 35787 29000 35829 29009
rect 35787 28960 35788 29000
rect 35828 28960 35829 29000
rect 35787 28951 35829 28960
rect 35788 28866 35828 28951
rect 35884 27077 35924 29044
rect 35883 27068 35925 27077
rect 35883 27028 35884 27068
rect 35924 27028 35925 27068
rect 35883 27019 35925 27028
rect 35596 26860 35732 26900
rect 34924 26767 34964 26776
rect 35308 26816 35348 26825
rect 34592 26480 34960 26489
rect 34632 26440 34674 26480
rect 34714 26440 34756 26480
rect 34796 26440 34838 26480
rect 34878 26440 34920 26480
rect 34592 26431 34960 26440
rect 34348 26095 34388 26104
rect 35308 26144 35348 26776
rect 35403 26816 35445 26825
rect 35403 26776 35404 26816
rect 35444 26776 35445 26816
rect 35403 26767 35445 26776
rect 35308 26069 35348 26104
rect 35307 26060 35349 26069
rect 35307 26020 35308 26060
rect 35348 26020 35349 26060
rect 35307 26011 35349 26020
rect 33352 25724 33720 25733
rect 33392 25684 33434 25724
rect 33474 25684 33516 25724
rect 33556 25684 33598 25724
rect 33638 25684 33680 25724
rect 33352 25675 33720 25684
rect 35211 25220 35253 25229
rect 35211 25180 35212 25220
rect 35252 25180 35253 25220
rect 35211 25171 35253 25180
rect 34592 24968 34960 24977
rect 34632 24928 34674 24968
rect 34714 24928 34756 24968
rect 34796 24928 34838 24968
rect 34878 24928 34920 24968
rect 34592 24919 34960 24928
rect 35212 24557 35252 25171
rect 35211 24548 35253 24557
rect 35211 24508 35212 24548
rect 35252 24508 35253 24548
rect 35211 24499 35253 24508
rect 33352 24212 33720 24221
rect 33392 24172 33434 24212
rect 33474 24172 33516 24212
rect 33556 24172 33598 24212
rect 33638 24172 33680 24212
rect 33352 24163 33720 24172
rect 32811 23876 32853 23885
rect 32811 23836 32812 23876
rect 32852 23836 32853 23876
rect 32811 23827 32853 23836
rect 30123 23792 30165 23801
rect 30123 23752 30124 23792
rect 30164 23752 30165 23792
rect 30123 23743 30165 23752
rect 29643 23708 29685 23717
rect 29643 23668 29644 23708
rect 29684 23668 29685 23708
rect 29643 23659 29685 23668
rect 32812 23633 32852 23827
rect 33292 23792 33332 23801
rect 33196 23752 33292 23792
rect 32811 23624 32853 23633
rect 32811 23584 32812 23624
rect 32852 23584 32853 23624
rect 32811 23575 32853 23584
rect 32619 22532 32661 22541
rect 32619 22492 32620 22532
rect 32660 22492 32661 22532
rect 32619 22483 32661 22492
rect 29163 20936 29205 20945
rect 29068 20896 29164 20936
rect 29204 20896 29205 20936
rect 29163 20887 29205 20896
rect 28875 20852 28917 20861
rect 28875 20812 28876 20852
rect 28916 20812 28917 20852
rect 28875 20803 28917 20812
rect 29164 20768 29204 20887
rect 29260 20777 29300 22240
rect 32428 22280 32468 22289
rect 32428 22121 32468 22240
rect 32523 22280 32565 22289
rect 32523 22240 32524 22280
rect 32564 22240 32565 22280
rect 32523 22231 32565 22240
rect 32620 22280 32660 22483
rect 32620 22231 32660 22240
rect 32524 22146 32564 22231
rect 32427 22112 32469 22121
rect 32427 22072 32428 22112
rect 32468 22072 32469 22112
rect 32427 22063 32469 22072
rect 33099 21860 33141 21869
rect 33099 21820 33100 21860
rect 33140 21820 33141 21860
rect 33099 21811 33141 21820
rect 29355 21608 29397 21617
rect 29355 21568 29356 21608
rect 29396 21568 29397 21608
rect 29355 21559 29397 21568
rect 29356 21474 29396 21559
rect 30315 20936 30357 20945
rect 30315 20896 30316 20936
rect 30356 20896 30357 20936
rect 30315 20887 30357 20896
rect 30604 20936 30644 20945
rect 30644 20896 30836 20936
rect 30604 20887 30644 20896
rect 29164 20719 29204 20728
rect 29259 20768 29301 20777
rect 29259 20728 29260 20768
rect 29300 20728 29301 20768
rect 29259 20719 29301 20728
rect 29643 20768 29685 20777
rect 29643 20728 29644 20768
rect 29684 20728 29685 20768
rect 29643 20719 29685 20728
rect 30316 20768 30356 20887
rect 30796 20852 30836 20896
rect 30796 20803 30836 20812
rect 31371 20852 31413 20861
rect 31371 20812 31372 20852
rect 31412 20812 31413 20852
rect 31371 20803 31413 20812
rect 30316 20719 30356 20728
rect 30507 20768 30549 20777
rect 30507 20728 30508 20768
rect 30548 20728 30549 20768
rect 30507 20719 30549 20728
rect 30604 20768 30644 20777
rect 29452 20600 29492 20609
rect 29452 20189 29492 20560
rect 29644 20600 29684 20719
rect 30508 20634 30548 20719
rect 29644 20551 29684 20560
rect 28107 20180 28149 20189
rect 28107 20140 28108 20180
rect 28148 20140 28149 20180
rect 28107 20131 28149 20140
rect 29451 20180 29493 20189
rect 29451 20140 29452 20180
rect 29492 20140 29493 20180
rect 29451 20131 29493 20140
rect 27339 18668 27381 18677
rect 27339 18628 27340 18668
rect 27380 18628 27381 18668
rect 27339 18619 27381 18628
rect 27340 18534 27380 18619
rect 27435 18584 27477 18593
rect 27435 18544 27436 18584
rect 27476 18544 27477 18584
rect 27435 18535 27477 18544
rect 27436 18450 27476 18535
rect 27148 17744 27188 17753
rect 27148 16997 27188 17704
rect 28011 17744 28053 17753
rect 28011 17704 28012 17744
rect 28052 17704 28053 17744
rect 28011 17695 28053 17704
rect 28012 17610 28052 17695
rect 28108 17492 28148 20131
rect 28395 18584 28437 18593
rect 28395 18544 28396 18584
rect 28436 18544 28437 18584
rect 28395 18535 28437 18544
rect 29068 18584 29108 18593
rect 29108 18544 29204 18584
rect 29068 18535 29108 18544
rect 28396 18450 28436 18535
rect 29164 17828 29204 18544
rect 29164 17669 29204 17788
rect 28203 17660 28245 17669
rect 28203 17620 28204 17660
rect 28244 17620 28245 17660
rect 28203 17611 28245 17620
rect 29163 17660 29205 17669
rect 29163 17620 29164 17660
rect 29204 17620 29205 17660
rect 29163 17611 29205 17620
rect 28012 17452 28148 17492
rect 27147 16988 27189 16997
rect 27147 16948 27148 16988
rect 27188 16948 27189 16988
rect 27147 16939 27189 16948
rect 27915 15560 27957 15569
rect 27915 15520 27916 15560
rect 27956 15520 27957 15560
rect 27915 15511 27957 15520
rect 27916 15426 27956 15511
rect 28012 15476 28052 17452
rect 28012 15427 28052 15436
rect 28204 15476 28244 17611
rect 30604 16409 30644 20728
rect 31180 20768 31220 20777
rect 30891 20600 30933 20609
rect 30891 20560 30892 20600
rect 30932 20560 30933 20600
rect 30891 20551 30933 20560
rect 30892 20466 30932 20551
rect 31180 16997 31220 20728
rect 31372 20718 31412 20803
rect 32619 18920 32661 18929
rect 32619 18880 32620 18920
rect 32660 18880 32661 18920
rect 32619 18871 32661 18880
rect 31371 17828 31413 17837
rect 31371 17788 31372 17828
rect 31412 17788 31413 17828
rect 31371 17779 31413 17788
rect 31372 17156 31412 17779
rect 32620 17753 32660 18871
rect 33100 17753 33140 21811
rect 33196 21617 33236 23752
rect 33292 23743 33332 23752
rect 34443 23792 34485 23801
rect 34443 23752 34444 23792
rect 34484 23752 34485 23792
rect 34443 23743 34485 23752
rect 33771 23624 33813 23633
rect 33771 23584 33772 23624
rect 33812 23584 33813 23624
rect 33771 23575 33813 23584
rect 33772 23490 33812 23575
rect 34060 23120 34100 23129
rect 33352 22700 33720 22709
rect 33392 22660 33434 22700
rect 33474 22660 33516 22700
rect 33556 22660 33598 22700
rect 33638 22660 33680 22700
rect 33352 22651 33720 22660
rect 34060 22448 34100 23080
rect 34444 23120 34484 23743
rect 34592 23456 34960 23465
rect 34632 23416 34674 23456
rect 34714 23416 34756 23456
rect 34796 23416 34838 23456
rect 34878 23416 34920 23456
rect 34592 23407 34960 23416
rect 34444 23071 34484 23080
rect 34155 22616 34197 22625
rect 34155 22576 34156 22616
rect 34196 22576 34197 22616
rect 34155 22567 34197 22576
rect 34923 22616 34965 22625
rect 34923 22576 34924 22616
rect 34964 22576 34965 22616
rect 34923 22567 34965 22576
rect 33964 22408 34100 22448
rect 33964 22028 34004 22408
rect 34059 22280 34101 22289
rect 34059 22240 34060 22280
rect 34100 22240 34101 22280
rect 34059 22231 34101 22240
rect 34156 22280 34196 22567
rect 34347 22364 34389 22373
rect 34347 22324 34348 22364
rect 34388 22324 34389 22364
rect 34347 22315 34389 22324
rect 34731 22364 34773 22373
rect 34731 22324 34732 22364
rect 34772 22324 34773 22364
rect 34731 22315 34773 22324
rect 34156 22231 34196 22240
rect 34060 22146 34100 22231
rect 34251 22196 34293 22205
rect 34251 22156 34252 22196
rect 34292 22156 34293 22196
rect 34251 22147 34293 22156
rect 34155 22112 34197 22121
rect 34155 22072 34156 22112
rect 34196 22072 34197 22112
rect 34155 22063 34197 22072
rect 33964 21988 34100 22028
rect 33195 21608 33237 21617
rect 33195 21568 33196 21608
rect 33236 21568 33237 21608
rect 33195 21559 33237 21568
rect 33196 19256 33236 21559
rect 33352 21188 33720 21197
rect 33392 21148 33434 21188
rect 33474 21148 33516 21188
rect 33556 21148 33598 21188
rect 33638 21148 33680 21188
rect 33352 21139 33720 21148
rect 34060 20693 34100 21988
rect 34059 20684 34101 20693
rect 34059 20644 34060 20684
rect 34100 20644 34101 20684
rect 34059 20635 34101 20644
rect 33771 20096 33813 20105
rect 33771 20056 33772 20096
rect 33812 20056 33813 20096
rect 33771 20047 33813 20056
rect 33352 19676 33720 19685
rect 33392 19636 33434 19676
rect 33474 19636 33516 19676
rect 33556 19636 33598 19676
rect 33638 19636 33680 19676
rect 33352 19627 33720 19636
rect 33196 19207 33236 19216
rect 33352 18164 33720 18173
rect 33392 18124 33434 18164
rect 33474 18124 33516 18164
rect 33556 18124 33598 18164
rect 33638 18124 33680 18164
rect 33352 18115 33720 18124
rect 33772 17996 33812 20047
rect 33868 19424 33908 19433
rect 33868 19265 33908 19384
rect 33867 19256 33909 19265
rect 33867 19216 33868 19256
rect 33908 19216 33909 19256
rect 33867 19207 33909 19216
rect 33868 18929 33908 19207
rect 33867 18920 33909 18929
rect 33867 18880 33868 18920
rect 33908 18880 33909 18920
rect 33867 18871 33909 18880
rect 33580 17956 33812 17996
rect 32619 17744 32661 17753
rect 32619 17704 32620 17744
rect 32660 17704 32661 17744
rect 32619 17695 32661 17704
rect 33099 17744 33141 17753
rect 33099 17704 33100 17744
rect 33140 17704 33141 17744
rect 33099 17695 33141 17704
rect 31372 17107 31412 17116
rect 31275 17072 31317 17081
rect 31275 17032 31276 17072
rect 31316 17032 31317 17072
rect 31275 17023 31317 17032
rect 31755 17072 31797 17081
rect 31755 17032 31756 17072
rect 31796 17032 31797 17072
rect 31755 17023 31797 17032
rect 32620 17072 32660 17695
rect 31179 16988 31221 16997
rect 31179 16948 31180 16988
rect 31220 16948 31221 16988
rect 31179 16939 31221 16948
rect 30603 16400 30645 16409
rect 30603 16360 30604 16400
rect 30644 16360 30645 16400
rect 30603 16351 30645 16360
rect 28300 15560 28340 15571
rect 28300 15485 28340 15520
rect 28204 15427 28244 15436
rect 28299 15476 28341 15485
rect 28299 15436 28300 15476
rect 28340 15436 28341 15476
rect 28299 15427 28341 15436
rect 28108 15392 28148 15401
rect 27819 12788 27861 12797
rect 27819 12748 27820 12788
rect 27860 12748 27861 12788
rect 27819 12739 27861 12748
rect 27243 12620 27285 12629
rect 27243 12580 27244 12620
rect 27284 12580 27285 12620
rect 27243 12571 27285 12580
rect 27244 12536 27284 12571
rect 27244 12485 27284 12496
rect 27820 12536 27860 12739
rect 27820 12487 27860 12496
rect 27435 12452 27477 12461
rect 27435 12412 27436 12452
rect 27476 12412 27477 12452
rect 27435 12403 27477 12412
rect 28011 12452 28053 12461
rect 28108 12452 28148 15352
rect 28011 12412 28012 12452
rect 28052 12412 28148 12452
rect 30892 12536 30932 12545
rect 28011 12403 28053 12412
rect 27436 12318 27476 12403
rect 28012 12318 28052 12403
rect 30700 12368 30740 12377
rect 30892 12368 30932 12496
rect 31276 12536 31316 17023
rect 31756 16938 31796 17023
rect 32620 15140 32660 17032
rect 33100 15569 33140 17695
rect 33580 16820 33620 17956
rect 33675 17744 33717 17753
rect 33675 17704 33676 17744
rect 33716 17704 33717 17744
rect 33675 17695 33717 17704
rect 33868 17744 33908 17753
rect 33676 17610 33716 17695
rect 33771 17660 33813 17669
rect 33771 17620 33772 17660
rect 33812 17620 33813 17660
rect 33771 17611 33813 17620
rect 33772 17526 33812 17611
rect 33772 16988 33812 16997
rect 33772 16904 33812 16948
rect 33868 16904 33908 17704
rect 34059 16988 34101 16997
rect 33772 16864 33908 16904
rect 33964 16948 34060 16988
rect 34100 16948 34101 16988
rect 33580 16780 33908 16820
rect 33352 16652 33720 16661
rect 33392 16612 33434 16652
rect 33474 16612 33516 16652
rect 33556 16612 33598 16652
rect 33638 16612 33680 16652
rect 33352 16603 33720 16612
rect 33195 16400 33237 16409
rect 33195 16360 33196 16400
rect 33236 16360 33237 16400
rect 33195 16351 33237 16360
rect 33771 16400 33813 16409
rect 33771 16360 33772 16400
rect 33812 16360 33813 16400
rect 33771 16351 33813 16360
rect 33099 15560 33141 15569
rect 33099 15520 33100 15560
rect 33140 15520 33141 15560
rect 33099 15511 33141 15520
rect 31276 12487 31316 12496
rect 32140 15100 32660 15140
rect 32140 12536 32180 15100
rect 33196 13460 33236 16351
rect 33772 16232 33812 16351
rect 33868 16316 33908 16780
rect 33964 16400 34004 16948
rect 34059 16939 34101 16948
rect 34060 16854 34100 16939
rect 33964 16351 34004 16360
rect 33868 16267 33908 16276
rect 34059 16316 34101 16325
rect 34059 16276 34060 16316
rect 34100 16276 34101 16316
rect 34059 16267 34101 16276
rect 33772 16183 33812 16192
rect 34060 16182 34100 16267
rect 34156 16232 34196 22063
rect 34252 22062 34292 22147
rect 34348 22112 34388 22315
rect 34636 22121 34676 22206
rect 34348 22063 34388 22072
rect 34444 22112 34484 22121
rect 34347 21944 34389 21953
rect 34347 21904 34348 21944
rect 34388 21904 34389 21944
rect 34347 21895 34389 21904
rect 34251 17660 34293 17669
rect 34251 17620 34252 17660
rect 34292 17620 34293 17660
rect 34251 17611 34293 17620
rect 34252 17072 34292 17611
rect 34252 17023 34292 17032
rect 33352 15140 33720 15149
rect 33392 15100 33434 15140
rect 33474 15100 33516 15140
rect 33556 15100 33598 15140
rect 33638 15100 33680 15140
rect 33352 15091 33720 15100
rect 33352 13628 33720 13637
rect 33392 13588 33434 13628
rect 33474 13588 33516 13628
rect 33556 13588 33598 13628
rect 33638 13588 33680 13628
rect 33352 13579 33720 13588
rect 33196 13420 33332 13460
rect 33195 13208 33237 13217
rect 33195 13168 33196 13208
rect 33236 13168 33237 13208
rect 33195 13159 33237 13168
rect 33196 13074 33236 13159
rect 33003 13040 33045 13049
rect 33003 13000 33004 13040
rect 33044 13000 33045 13040
rect 33003 12991 33045 13000
rect 33292 13040 33332 13420
rect 34156 13217 34196 16192
rect 34252 16820 34292 16829
rect 34155 13208 34197 13217
rect 34155 13168 34156 13208
rect 34196 13168 34197 13208
rect 34155 13159 34197 13168
rect 33004 12906 33044 12991
rect 32140 12487 32180 12496
rect 33292 12536 33332 13000
rect 33292 12487 33332 12496
rect 30740 12328 30932 12368
rect 30700 12319 30740 12328
rect 27243 12284 27285 12293
rect 27243 12244 27244 12284
rect 27284 12244 27285 12284
rect 27243 12235 27285 12244
rect 27820 12284 27860 12293
rect 27244 12150 27284 12235
rect 27820 12041 27860 12244
rect 33352 12116 33720 12125
rect 33392 12076 33434 12116
rect 33474 12076 33516 12116
rect 33556 12076 33598 12116
rect 33638 12076 33680 12116
rect 33352 12067 33720 12076
rect 27819 12032 27861 12041
rect 27819 11992 27820 12032
rect 27860 11992 27861 12032
rect 27819 11983 27861 11992
rect 33352 10604 33720 10613
rect 33392 10564 33434 10604
rect 33474 10564 33516 10604
rect 33556 10564 33598 10604
rect 33638 10564 33680 10604
rect 33352 10555 33720 10564
rect 27051 9428 27093 9437
rect 27051 9388 27052 9428
rect 27092 9388 27093 9428
rect 27051 9379 27093 9388
rect 33352 9092 33720 9101
rect 33392 9052 33434 9092
rect 33474 9052 33516 9092
rect 33556 9052 33598 9092
rect 33638 9052 33680 9092
rect 33352 9043 33720 9052
rect 19472 8336 19840 8345
rect 19512 8296 19554 8336
rect 19594 8296 19636 8336
rect 19676 8296 19718 8336
rect 19758 8296 19800 8336
rect 19472 8287 19840 8296
rect 33352 7580 33720 7589
rect 33392 7540 33434 7580
rect 33474 7540 33516 7580
rect 33556 7540 33598 7580
rect 33638 7540 33680 7580
rect 33352 7531 33720 7540
rect 34252 7253 34292 16780
rect 34251 7244 34293 7253
rect 34251 7204 34252 7244
rect 34292 7204 34293 7244
rect 34251 7195 34293 7204
rect 19472 6824 19840 6833
rect 19512 6784 19554 6824
rect 19594 6784 19636 6824
rect 19676 6784 19718 6824
rect 19758 6784 19800 6824
rect 19472 6775 19840 6784
rect 18700 6280 18836 6320
rect 3112 6068 3480 6077
rect 3152 6028 3194 6068
rect 3234 6028 3276 6068
rect 3316 6028 3358 6068
rect 3398 6028 3440 6068
rect 3112 6019 3480 6028
rect 18232 6068 18600 6077
rect 18272 6028 18314 6068
rect 18354 6028 18396 6068
rect 18436 6028 18478 6068
rect 18518 6028 18560 6068
rect 18232 6019 18600 6028
rect 18700 5741 18740 6280
rect 33352 6068 33720 6077
rect 33392 6028 33434 6068
rect 33474 6028 33516 6068
rect 33556 6028 33598 6068
rect 33638 6028 33680 6068
rect 33352 6019 33720 6028
rect 18699 5732 18741 5741
rect 18699 5692 18700 5732
rect 18740 5692 18741 5732
rect 18699 5683 18741 5692
rect 4352 5312 4720 5321
rect 4392 5272 4434 5312
rect 4474 5272 4516 5312
rect 4556 5272 4598 5312
rect 4638 5272 4680 5312
rect 4352 5263 4720 5272
rect 19472 5312 19840 5321
rect 19512 5272 19554 5312
rect 19594 5272 19636 5312
rect 19676 5272 19718 5312
rect 19758 5272 19800 5312
rect 19472 5263 19840 5272
rect 34348 4901 34388 21895
rect 34347 4892 34389 4901
rect 34347 4852 34348 4892
rect 34388 4852 34389 4892
rect 34347 4843 34389 4852
rect 3112 4556 3480 4565
rect 3152 4516 3194 4556
rect 3234 4516 3276 4556
rect 3316 4516 3358 4556
rect 3398 4516 3440 4556
rect 3112 4507 3480 4516
rect 18232 4556 18600 4565
rect 18272 4516 18314 4556
rect 18354 4516 18396 4556
rect 18436 4516 18478 4556
rect 18518 4516 18560 4556
rect 18232 4507 18600 4516
rect 33352 4556 33720 4565
rect 33392 4516 33434 4556
rect 33474 4516 33516 4556
rect 33556 4516 33598 4556
rect 33638 4516 33680 4556
rect 33352 4507 33720 4516
rect 34444 4229 34484 22072
rect 34635 22112 34677 22121
rect 34635 22072 34636 22112
rect 34676 22072 34677 22112
rect 34635 22063 34677 22072
rect 34732 22112 34772 22315
rect 34924 22280 34964 22567
rect 34924 22231 34964 22240
rect 35020 22280 35060 22291
rect 35020 22205 35060 22240
rect 35212 22280 35252 24499
rect 35404 23633 35444 26767
rect 35499 26060 35541 26069
rect 35499 26020 35500 26060
rect 35540 26020 35541 26060
rect 35499 26011 35541 26020
rect 35500 23885 35540 26011
rect 35596 25229 35636 26860
rect 35595 25220 35637 25229
rect 35595 25180 35596 25220
rect 35636 25180 35637 25220
rect 35595 25171 35637 25180
rect 36076 23960 36116 29128
rect 36460 29009 36500 29800
rect 36748 29672 36788 29681
rect 36459 29000 36501 29009
rect 36459 28960 36460 29000
rect 36500 28960 36501 29000
rect 36459 28951 36501 28960
rect 36171 26816 36213 26825
rect 36171 26776 36172 26816
rect 36212 26776 36213 26816
rect 36171 26767 36213 26776
rect 36172 26682 36212 26767
rect 35980 23920 36116 23960
rect 35499 23876 35541 23885
rect 35499 23836 35500 23876
rect 35540 23836 35541 23876
rect 35499 23827 35541 23836
rect 35403 23624 35445 23633
rect 35403 23584 35404 23624
rect 35444 23584 35445 23624
rect 35403 23575 35445 23584
rect 35307 23120 35349 23129
rect 35404 23120 35444 23575
rect 35307 23080 35308 23120
rect 35348 23080 35444 23120
rect 35307 23071 35349 23080
rect 35308 22986 35348 23071
rect 35980 22457 36020 23920
rect 36460 22868 36500 22877
rect 35595 22448 35637 22457
rect 35595 22408 35596 22448
rect 35636 22408 35637 22448
rect 35595 22399 35637 22408
rect 35979 22448 36021 22457
rect 35979 22408 35980 22448
rect 36020 22408 36021 22448
rect 35979 22399 36021 22408
rect 35307 22364 35349 22373
rect 35307 22324 35308 22364
rect 35348 22324 35349 22364
rect 35307 22315 35349 22324
rect 34820 22196 34860 22205
rect 34820 22121 34860 22156
rect 35019 22196 35061 22205
rect 35019 22156 35020 22196
rect 35060 22156 35061 22196
rect 35019 22147 35061 22156
rect 34820 22112 34869 22121
rect 34820 22072 34828 22112
rect 34868 22072 34869 22112
rect 34732 22063 34772 22072
rect 34827 22063 34869 22072
rect 35019 22028 35061 22037
rect 35019 21988 35020 22028
rect 35060 21988 35061 22028
rect 35019 21979 35061 21988
rect 34592 21944 34960 21953
rect 34632 21904 34674 21944
rect 34714 21904 34756 21944
rect 34796 21904 34838 21944
rect 34878 21904 34920 21944
rect 34592 21895 34960 21904
rect 34592 20432 34960 20441
rect 34632 20392 34674 20432
rect 34714 20392 34756 20432
rect 34796 20392 34838 20432
rect 34878 20392 34920 20432
rect 34592 20383 34960 20392
rect 35020 20264 35060 21979
rect 35212 21869 35252 22240
rect 35308 22230 35348 22315
rect 35403 22280 35445 22289
rect 35403 22240 35404 22280
rect 35444 22240 35445 22280
rect 35403 22231 35445 22240
rect 35596 22280 35636 22399
rect 35787 22364 35829 22373
rect 35787 22324 35788 22364
rect 35828 22324 35829 22364
rect 35787 22315 35829 22324
rect 35596 22231 35636 22240
rect 35788 22280 35828 22315
rect 36460 22289 36500 22828
rect 35404 22146 35444 22231
rect 35788 22229 35828 22240
rect 36459 22280 36501 22289
rect 36459 22240 36460 22280
rect 36500 22240 36501 22280
rect 36459 22231 36501 22240
rect 35691 22196 35733 22205
rect 35691 22156 35692 22196
rect 35732 22156 35733 22196
rect 35691 22147 35733 22156
rect 35692 22062 35732 22147
rect 35211 21860 35253 21869
rect 35211 21820 35212 21860
rect 35252 21820 35253 21860
rect 35211 21811 35253 21820
rect 34924 20224 35060 20264
rect 34924 20180 34964 20224
rect 34924 20131 34964 20140
rect 34827 20096 34869 20105
rect 34827 20056 34828 20096
rect 34868 20056 34869 20096
rect 34827 20047 34869 20056
rect 35019 20096 35061 20105
rect 35019 20056 35020 20096
rect 35060 20056 35061 20096
rect 35019 20047 35061 20056
rect 34828 19962 34868 20047
rect 35020 19962 35060 20047
rect 34592 18920 34960 18929
rect 34632 18880 34674 18920
rect 34714 18880 34756 18920
rect 34796 18880 34838 18920
rect 34878 18880 34920 18920
rect 34592 18871 34960 18880
rect 34592 17408 34960 17417
rect 34632 17368 34674 17408
rect 34714 17368 34756 17408
rect 34796 17368 34838 17408
rect 34878 17368 34920 17408
rect 34592 17359 34960 17368
rect 34592 15896 34960 15905
rect 34632 15856 34674 15896
rect 34714 15856 34756 15896
rect 34796 15856 34838 15896
rect 34878 15856 34920 15896
rect 34592 15847 34960 15856
rect 34592 14384 34960 14393
rect 34632 14344 34674 14384
rect 34714 14344 34756 14384
rect 34796 14344 34838 14384
rect 34878 14344 34920 14384
rect 34592 14335 34960 14344
rect 34592 12872 34960 12881
rect 34632 12832 34674 12872
rect 34714 12832 34756 12872
rect 34796 12832 34838 12872
rect 34878 12832 34920 12872
rect 34592 12823 34960 12832
rect 34592 11360 34960 11369
rect 34632 11320 34674 11360
rect 34714 11320 34756 11360
rect 34796 11320 34838 11360
rect 34878 11320 34920 11360
rect 34592 11311 34960 11320
rect 36748 10277 36788 29632
rect 49712 29504 50080 29513
rect 49752 29464 49794 29504
rect 49834 29464 49876 29504
rect 49916 29464 49958 29504
rect 49998 29464 50040 29504
rect 49712 29455 50080 29464
rect 64832 29504 65200 29513
rect 64872 29464 64914 29504
rect 64954 29464 64996 29504
rect 65036 29464 65078 29504
rect 65118 29464 65160 29504
rect 64832 29455 65200 29464
rect 79952 29504 80320 29513
rect 79992 29464 80034 29504
rect 80074 29464 80116 29504
rect 80156 29464 80198 29504
rect 80238 29464 80280 29504
rect 79952 29455 80320 29464
rect 95072 29504 95440 29513
rect 95112 29464 95154 29504
rect 95194 29464 95236 29504
rect 95276 29464 95318 29504
rect 95358 29464 95400 29504
rect 95072 29455 95440 29464
rect 48472 28748 48840 28757
rect 48512 28708 48554 28748
rect 48594 28708 48636 28748
rect 48676 28708 48718 28748
rect 48758 28708 48800 28748
rect 48472 28699 48840 28708
rect 63592 28748 63960 28757
rect 63632 28708 63674 28748
rect 63714 28708 63756 28748
rect 63796 28708 63838 28748
rect 63878 28708 63920 28748
rect 63592 28699 63960 28708
rect 78712 28748 79080 28757
rect 78752 28708 78794 28748
rect 78834 28708 78876 28748
rect 78916 28708 78958 28748
rect 78998 28708 79040 28748
rect 78712 28699 79080 28708
rect 93832 28748 94200 28757
rect 93872 28708 93914 28748
rect 93954 28708 93996 28748
rect 94036 28708 94078 28748
rect 94118 28708 94160 28748
rect 93832 28699 94200 28708
rect 49712 27992 50080 28001
rect 49752 27952 49794 27992
rect 49834 27952 49876 27992
rect 49916 27952 49958 27992
rect 49998 27952 50040 27992
rect 49712 27943 50080 27952
rect 64832 27992 65200 28001
rect 64872 27952 64914 27992
rect 64954 27952 64996 27992
rect 65036 27952 65078 27992
rect 65118 27952 65160 27992
rect 64832 27943 65200 27952
rect 79952 27992 80320 28001
rect 79992 27952 80034 27992
rect 80074 27952 80116 27992
rect 80156 27952 80198 27992
rect 80238 27952 80280 27992
rect 79952 27943 80320 27952
rect 95072 27992 95440 28001
rect 95112 27952 95154 27992
rect 95194 27952 95236 27992
rect 95276 27952 95318 27992
rect 95358 27952 95400 27992
rect 95072 27943 95440 27952
rect 48472 27236 48840 27245
rect 48512 27196 48554 27236
rect 48594 27196 48636 27236
rect 48676 27196 48718 27236
rect 48758 27196 48800 27236
rect 48472 27187 48840 27196
rect 63592 27236 63960 27245
rect 63632 27196 63674 27236
rect 63714 27196 63756 27236
rect 63796 27196 63838 27236
rect 63878 27196 63920 27236
rect 63592 27187 63960 27196
rect 78712 27236 79080 27245
rect 78752 27196 78794 27236
rect 78834 27196 78876 27236
rect 78916 27196 78958 27236
rect 78998 27196 79040 27236
rect 78712 27187 79080 27196
rect 93832 27236 94200 27245
rect 93872 27196 93914 27236
rect 93954 27196 93996 27236
rect 94036 27196 94078 27236
rect 94118 27196 94160 27236
rect 93832 27187 94200 27196
rect 37323 27068 37365 27077
rect 37323 27028 37324 27068
rect 37364 27028 37365 27068
rect 37323 27019 37365 27028
rect 37324 26934 37364 27019
rect 49712 26480 50080 26489
rect 49752 26440 49794 26480
rect 49834 26440 49876 26480
rect 49916 26440 49958 26480
rect 49998 26440 50040 26480
rect 49712 26431 50080 26440
rect 64832 26480 65200 26489
rect 64872 26440 64914 26480
rect 64954 26440 64996 26480
rect 65036 26440 65078 26480
rect 65118 26440 65160 26480
rect 64832 26431 65200 26440
rect 79952 26480 80320 26489
rect 79992 26440 80034 26480
rect 80074 26440 80116 26480
rect 80156 26440 80198 26480
rect 80238 26440 80280 26480
rect 79952 26431 80320 26440
rect 95072 26480 95440 26489
rect 95112 26440 95154 26480
rect 95194 26440 95236 26480
rect 95276 26440 95318 26480
rect 95358 26440 95400 26480
rect 95072 26431 95440 26440
rect 39627 26144 39669 26153
rect 39627 26104 39628 26144
rect 39668 26104 39669 26144
rect 39627 26095 39669 26104
rect 39628 26010 39668 26095
rect 39916 25892 39956 25901
rect 39916 23885 39956 25852
rect 48472 25724 48840 25733
rect 48512 25684 48554 25724
rect 48594 25684 48636 25724
rect 48676 25684 48718 25724
rect 48758 25684 48800 25724
rect 48472 25675 48840 25684
rect 63592 25724 63960 25733
rect 63632 25684 63674 25724
rect 63714 25684 63756 25724
rect 63796 25684 63838 25724
rect 63878 25684 63920 25724
rect 63592 25675 63960 25684
rect 78712 25724 79080 25733
rect 78752 25684 78794 25724
rect 78834 25684 78876 25724
rect 78916 25684 78958 25724
rect 78998 25684 79040 25724
rect 78712 25675 79080 25684
rect 93832 25724 94200 25733
rect 93872 25684 93914 25724
rect 93954 25684 93996 25724
rect 94036 25684 94078 25724
rect 94118 25684 94160 25724
rect 93832 25675 94200 25684
rect 49712 24968 50080 24977
rect 49752 24928 49794 24968
rect 49834 24928 49876 24968
rect 49916 24928 49958 24968
rect 49998 24928 50040 24968
rect 49712 24919 50080 24928
rect 64832 24968 65200 24977
rect 64872 24928 64914 24968
rect 64954 24928 64996 24968
rect 65036 24928 65078 24968
rect 65118 24928 65160 24968
rect 64832 24919 65200 24928
rect 79952 24968 80320 24977
rect 79992 24928 80034 24968
rect 80074 24928 80116 24968
rect 80156 24928 80198 24968
rect 80238 24928 80280 24968
rect 79952 24919 80320 24928
rect 95072 24968 95440 24977
rect 95112 24928 95154 24968
rect 95194 24928 95236 24968
rect 95276 24928 95318 24968
rect 95358 24928 95400 24968
rect 95072 24919 95440 24928
rect 48472 24212 48840 24221
rect 48512 24172 48554 24212
rect 48594 24172 48636 24212
rect 48676 24172 48718 24212
rect 48758 24172 48800 24212
rect 48472 24163 48840 24172
rect 63592 24212 63960 24221
rect 63632 24172 63674 24212
rect 63714 24172 63756 24212
rect 63796 24172 63838 24212
rect 63878 24172 63920 24212
rect 63592 24163 63960 24172
rect 78712 24212 79080 24221
rect 78752 24172 78794 24212
rect 78834 24172 78876 24212
rect 78916 24172 78958 24212
rect 78998 24172 79040 24212
rect 78712 24163 79080 24172
rect 93832 24212 94200 24221
rect 93872 24172 93914 24212
rect 93954 24172 93996 24212
rect 94036 24172 94078 24212
rect 94118 24172 94160 24212
rect 93832 24163 94200 24172
rect 39915 23876 39957 23885
rect 39915 23836 39916 23876
rect 39956 23836 39957 23876
rect 39915 23827 39957 23836
rect 39916 22709 39956 23827
rect 49712 23456 50080 23465
rect 49752 23416 49794 23456
rect 49834 23416 49876 23456
rect 49916 23416 49958 23456
rect 49998 23416 50040 23456
rect 49712 23407 50080 23416
rect 64832 23456 65200 23465
rect 64872 23416 64914 23456
rect 64954 23416 64996 23456
rect 65036 23416 65078 23456
rect 65118 23416 65160 23456
rect 64832 23407 65200 23416
rect 79952 23456 80320 23465
rect 79992 23416 80034 23456
rect 80074 23416 80116 23456
rect 80156 23416 80198 23456
rect 80238 23416 80280 23456
rect 79952 23407 80320 23416
rect 95072 23456 95440 23465
rect 95112 23416 95154 23456
rect 95194 23416 95236 23456
rect 95276 23416 95318 23456
rect 95358 23416 95400 23456
rect 95072 23407 95440 23416
rect 40395 23120 40437 23129
rect 40395 23080 40396 23120
rect 40436 23080 40437 23120
rect 40395 23071 40437 23080
rect 39531 22700 39573 22709
rect 39531 22660 39532 22700
rect 39572 22660 39573 22700
rect 39531 22651 39573 22660
rect 39915 22700 39957 22709
rect 39915 22660 39916 22700
rect 39956 22660 39957 22700
rect 39915 22651 39957 22660
rect 39532 22280 39572 22651
rect 39148 22196 39188 22205
rect 39052 22156 39148 22196
rect 37227 19844 37269 19853
rect 37227 19804 37228 19844
rect 37268 19804 37269 19844
rect 37227 19795 37269 19804
rect 37035 19340 37077 19349
rect 37035 19300 37036 19340
rect 37076 19300 37172 19340
rect 37035 19291 37077 19300
rect 36844 19256 36884 19265
rect 36844 18677 36884 19216
rect 37132 19256 37172 19300
rect 37132 19207 37172 19216
rect 37228 19256 37268 19795
rect 37515 19424 37557 19433
rect 37515 19384 37516 19424
rect 37556 19384 37557 19424
rect 37515 19375 37557 19384
rect 38763 19424 38805 19433
rect 38763 19384 38764 19424
rect 38804 19384 38805 19424
rect 38763 19375 38805 19384
rect 37516 19290 37556 19375
rect 37228 19207 37268 19216
rect 38764 19256 38804 19375
rect 38764 19207 38804 19216
rect 38859 19256 38901 19265
rect 38859 19216 38860 19256
rect 38900 19216 38901 19256
rect 38859 19207 38901 19216
rect 38763 19088 38805 19097
rect 38763 19048 38764 19088
rect 38804 19048 38805 19088
rect 38763 19039 38805 19048
rect 36843 18668 36885 18677
rect 36843 18628 36844 18668
rect 36884 18628 36885 18668
rect 36843 18619 36885 18628
rect 37227 18668 37269 18677
rect 37227 18628 37228 18668
rect 37268 18628 37269 18668
rect 37227 18619 37269 18628
rect 37228 16232 37268 18619
rect 37900 17744 37940 17753
rect 37900 17165 37940 17704
rect 38764 17744 38804 19039
rect 38764 17695 38804 17704
rect 37899 17156 37941 17165
rect 37899 17116 37900 17156
rect 37940 17116 37941 17156
rect 37899 17107 37941 17116
rect 37228 16183 37268 16192
rect 37323 16232 37365 16241
rect 37323 16192 37324 16232
rect 37364 16192 37365 16232
rect 37323 16183 37365 16192
rect 37324 16098 37364 16183
rect 37036 16064 37076 16073
rect 37036 15644 37076 16024
rect 37612 15644 37652 15653
rect 37036 15604 37612 15644
rect 37612 15595 37652 15604
rect 37900 15560 37940 17107
rect 38571 16232 38613 16241
rect 38571 16192 38572 16232
rect 38612 16192 38613 16232
rect 38571 16183 38613 16192
rect 38572 16098 38612 16183
rect 37996 15560 38036 15569
rect 37900 15520 37996 15560
rect 37996 15511 38036 15520
rect 38860 15560 38900 19207
rect 39052 18509 39092 22156
rect 39148 22147 39188 22156
rect 39243 19844 39285 19853
rect 39243 19804 39244 19844
rect 39284 19804 39285 19844
rect 39243 19795 39285 19804
rect 39244 19710 39284 19795
rect 39148 19256 39188 19265
rect 39148 19097 39188 19216
rect 39532 19097 39572 22240
rect 40396 22280 40436 23071
rect 48472 22700 48840 22709
rect 48512 22660 48554 22700
rect 48594 22660 48636 22700
rect 48676 22660 48718 22700
rect 48758 22660 48800 22700
rect 48472 22651 48840 22660
rect 63592 22700 63960 22709
rect 63632 22660 63674 22700
rect 63714 22660 63756 22700
rect 63796 22660 63838 22700
rect 63878 22660 63920 22700
rect 63592 22651 63960 22660
rect 78712 22700 79080 22709
rect 78752 22660 78794 22700
rect 78834 22660 78876 22700
rect 78916 22660 78958 22700
rect 78998 22660 79040 22700
rect 78712 22651 79080 22660
rect 93832 22700 94200 22709
rect 93872 22660 93914 22700
rect 93954 22660 93996 22700
rect 94036 22660 94078 22700
rect 94118 22660 94160 22700
rect 93832 22651 94200 22660
rect 41547 22364 41589 22373
rect 41547 22324 41548 22364
rect 41588 22324 41589 22364
rect 41547 22315 41589 22324
rect 40396 22231 40436 22240
rect 41548 22230 41588 22315
rect 49712 21944 50080 21953
rect 49752 21904 49794 21944
rect 49834 21904 49876 21944
rect 49916 21904 49958 21944
rect 49998 21904 50040 21944
rect 49712 21895 50080 21904
rect 64832 21944 65200 21953
rect 64872 21904 64914 21944
rect 64954 21904 64996 21944
rect 65036 21904 65078 21944
rect 65118 21904 65160 21944
rect 64832 21895 65200 21904
rect 79952 21944 80320 21953
rect 79992 21904 80034 21944
rect 80074 21904 80116 21944
rect 80156 21904 80198 21944
rect 80238 21904 80280 21944
rect 79952 21895 80320 21904
rect 95072 21944 95440 21953
rect 95112 21904 95154 21944
rect 95194 21904 95236 21944
rect 95276 21904 95318 21944
rect 95358 21904 95400 21944
rect 95072 21895 95440 21904
rect 48472 21188 48840 21197
rect 48512 21148 48554 21188
rect 48594 21148 48636 21188
rect 48676 21148 48718 21188
rect 48758 21148 48800 21188
rect 48472 21139 48840 21148
rect 63592 21188 63960 21197
rect 63632 21148 63674 21188
rect 63714 21148 63756 21188
rect 63796 21148 63838 21188
rect 63878 21148 63920 21188
rect 63592 21139 63960 21148
rect 78712 21188 79080 21197
rect 78752 21148 78794 21188
rect 78834 21148 78876 21188
rect 78916 21148 78958 21188
rect 78998 21148 79040 21188
rect 78712 21139 79080 21148
rect 93832 21188 94200 21197
rect 93872 21148 93914 21188
rect 93954 21148 93996 21188
rect 94036 21148 94078 21188
rect 94118 21148 94160 21188
rect 93832 21139 94200 21148
rect 49712 20432 50080 20441
rect 49752 20392 49794 20432
rect 49834 20392 49876 20432
rect 49916 20392 49958 20432
rect 49998 20392 50040 20432
rect 49712 20383 50080 20392
rect 64832 20432 65200 20441
rect 64872 20392 64914 20432
rect 64954 20392 64996 20432
rect 65036 20392 65078 20432
rect 65118 20392 65160 20432
rect 64832 20383 65200 20392
rect 79952 20432 80320 20441
rect 79992 20392 80034 20432
rect 80074 20392 80116 20432
rect 80156 20392 80198 20432
rect 80238 20392 80280 20432
rect 79952 20383 80320 20392
rect 95072 20432 95440 20441
rect 95112 20392 95154 20432
rect 95194 20392 95236 20432
rect 95276 20392 95318 20432
rect 95358 20392 95400 20432
rect 95072 20383 95440 20392
rect 39915 20096 39957 20105
rect 39915 20056 39916 20096
rect 39956 20056 39957 20096
rect 39915 20047 39957 20056
rect 41163 20096 41205 20105
rect 41163 20056 41164 20096
rect 41204 20056 41205 20096
rect 41163 20047 41205 20056
rect 39916 19962 39956 20047
rect 41164 19508 41204 20047
rect 48472 19676 48840 19685
rect 48512 19636 48554 19676
rect 48594 19636 48636 19676
rect 48676 19636 48718 19676
rect 48758 19636 48800 19676
rect 48472 19627 48840 19636
rect 63592 19676 63960 19685
rect 63632 19636 63674 19676
rect 63714 19636 63756 19676
rect 63796 19636 63838 19676
rect 63878 19636 63920 19676
rect 63592 19627 63960 19636
rect 78712 19676 79080 19685
rect 78752 19636 78794 19676
rect 78834 19636 78876 19676
rect 78916 19636 78958 19676
rect 78998 19636 79040 19676
rect 78712 19627 79080 19636
rect 93832 19676 94200 19685
rect 93872 19636 93914 19676
rect 93954 19636 93996 19676
rect 94036 19636 94078 19676
rect 94118 19636 94160 19676
rect 93832 19627 94200 19636
rect 41164 19459 41204 19468
rect 40011 19256 40053 19265
rect 40011 19216 40012 19256
rect 40052 19216 40053 19256
rect 40011 19207 40053 19216
rect 40012 19122 40052 19207
rect 39147 19088 39189 19097
rect 39147 19048 39148 19088
rect 39188 19048 39189 19088
rect 39147 19039 39189 19048
rect 39531 19088 39573 19097
rect 39531 19048 39532 19088
rect 39572 19048 39573 19088
rect 39531 19039 39573 19048
rect 49712 18920 50080 18929
rect 49752 18880 49794 18920
rect 49834 18880 49876 18920
rect 49916 18880 49958 18920
rect 49998 18880 50040 18920
rect 49712 18871 50080 18880
rect 64832 18920 65200 18929
rect 64872 18880 64914 18920
rect 64954 18880 64996 18920
rect 65036 18880 65078 18920
rect 65118 18880 65160 18920
rect 64832 18871 65200 18880
rect 79952 18920 80320 18929
rect 79992 18880 80034 18920
rect 80074 18880 80116 18920
rect 80156 18880 80198 18920
rect 80238 18880 80280 18920
rect 79952 18871 80320 18880
rect 95072 18920 95440 18929
rect 95112 18880 95154 18920
rect 95194 18880 95236 18920
rect 95276 18880 95318 18920
rect 95358 18880 95400 18920
rect 95072 18871 95440 18880
rect 39051 18500 39093 18509
rect 39051 18460 39052 18500
rect 39092 18460 39093 18500
rect 39051 18451 39093 18460
rect 48472 18164 48840 18173
rect 48512 18124 48554 18164
rect 48594 18124 48636 18164
rect 48676 18124 48718 18164
rect 48758 18124 48800 18164
rect 48472 18115 48840 18124
rect 63592 18164 63960 18173
rect 63632 18124 63674 18164
rect 63714 18124 63756 18164
rect 63796 18124 63838 18164
rect 63878 18124 63920 18164
rect 63592 18115 63960 18124
rect 78712 18164 79080 18173
rect 78752 18124 78794 18164
rect 78834 18124 78876 18164
rect 78916 18124 78958 18164
rect 78998 18124 79040 18164
rect 78712 18115 79080 18124
rect 93832 18164 94200 18173
rect 93872 18124 93914 18164
rect 93954 18124 93996 18164
rect 94036 18124 94078 18164
rect 94118 18124 94160 18164
rect 93832 18115 94200 18124
rect 49712 17408 50080 17417
rect 49752 17368 49794 17408
rect 49834 17368 49876 17408
rect 49916 17368 49958 17408
rect 49998 17368 50040 17408
rect 49712 17359 50080 17368
rect 64832 17408 65200 17417
rect 64872 17368 64914 17408
rect 64954 17368 64996 17408
rect 65036 17368 65078 17408
rect 65118 17368 65160 17408
rect 64832 17359 65200 17368
rect 79952 17408 80320 17417
rect 79992 17368 80034 17408
rect 80074 17368 80116 17408
rect 80156 17368 80198 17408
rect 80238 17368 80280 17408
rect 79952 17359 80320 17368
rect 95072 17408 95440 17417
rect 95112 17368 95154 17408
rect 95194 17368 95236 17408
rect 95276 17368 95318 17408
rect 95358 17368 95400 17408
rect 95072 17359 95440 17368
rect 48472 16652 48840 16661
rect 48512 16612 48554 16652
rect 48594 16612 48636 16652
rect 48676 16612 48718 16652
rect 48758 16612 48800 16652
rect 48472 16603 48840 16612
rect 63592 16652 63960 16661
rect 63632 16612 63674 16652
rect 63714 16612 63756 16652
rect 63796 16612 63838 16652
rect 63878 16612 63920 16652
rect 63592 16603 63960 16612
rect 78712 16652 79080 16661
rect 78752 16612 78794 16652
rect 78834 16612 78876 16652
rect 78916 16612 78958 16652
rect 78998 16612 79040 16652
rect 78712 16603 79080 16612
rect 93832 16652 94200 16661
rect 93872 16612 93914 16652
rect 93954 16612 93996 16652
rect 94036 16612 94078 16652
rect 94118 16612 94160 16652
rect 93832 16603 94200 16612
rect 39243 16316 39285 16325
rect 39243 16276 39244 16316
rect 39284 16276 39285 16316
rect 39243 16267 39285 16276
rect 40011 16316 40053 16325
rect 40011 16276 40012 16316
rect 40052 16276 40053 16316
rect 40011 16267 40053 16276
rect 39244 16232 39284 16267
rect 39244 16181 39284 16192
rect 40012 15728 40052 16267
rect 49712 15896 50080 15905
rect 49752 15856 49794 15896
rect 49834 15856 49876 15896
rect 49916 15856 49958 15896
rect 49998 15856 50040 15896
rect 49712 15847 50080 15856
rect 64832 15896 65200 15905
rect 64872 15856 64914 15896
rect 64954 15856 64996 15896
rect 65036 15856 65078 15896
rect 65118 15856 65160 15896
rect 64832 15847 65200 15856
rect 79952 15896 80320 15905
rect 79992 15856 80034 15896
rect 80074 15856 80116 15896
rect 80156 15856 80198 15896
rect 80238 15856 80280 15896
rect 79952 15847 80320 15856
rect 95072 15896 95440 15905
rect 95112 15856 95154 15896
rect 95194 15856 95236 15896
rect 95276 15856 95318 15896
rect 95358 15856 95400 15896
rect 95072 15847 95440 15856
rect 40012 15679 40052 15688
rect 38860 15511 38900 15520
rect 48472 15140 48840 15149
rect 48512 15100 48554 15140
rect 48594 15100 48636 15140
rect 48676 15100 48718 15140
rect 48758 15100 48800 15140
rect 48472 15091 48840 15100
rect 63592 15140 63960 15149
rect 63632 15100 63674 15140
rect 63714 15100 63756 15140
rect 63796 15100 63838 15140
rect 63878 15100 63920 15140
rect 63592 15091 63960 15100
rect 78712 15140 79080 15149
rect 78752 15100 78794 15140
rect 78834 15100 78876 15140
rect 78916 15100 78958 15140
rect 78998 15100 79040 15140
rect 78712 15091 79080 15100
rect 93832 15140 94200 15149
rect 93872 15100 93914 15140
rect 93954 15100 93996 15140
rect 94036 15100 94078 15140
rect 94118 15100 94160 15140
rect 93832 15091 94200 15100
rect 49712 14384 50080 14393
rect 49752 14344 49794 14384
rect 49834 14344 49876 14384
rect 49916 14344 49958 14384
rect 49998 14344 50040 14384
rect 49712 14335 50080 14344
rect 64832 14384 65200 14393
rect 64872 14344 64914 14384
rect 64954 14344 64996 14384
rect 65036 14344 65078 14384
rect 65118 14344 65160 14384
rect 64832 14335 65200 14344
rect 79952 14384 80320 14393
rect 79992 14344 80034 14384
rect 80074 14344 80116 14384
rect 80156 14344 80198 14384
rect 80238 14344 80280 14384
rect 79952 14335 80320 14344
rect 95072 14384 95440 14393
rect 95112 14344 95154 14384
rect 95194 14344 95236 14384
rect 95276 14344 95318 14384
rect 95358 14344 95400 14384
rect 95072 14335 95440 14344
rect 48472 13628 48840 13637
rect 48512 13588 48554 13628
rect 48594 13588 48636 13628
rect 48676 13588 48718 13628
rect 48758 13588 48800 13628
rect 48472 13579 48840 13588
rect 63592 13628 63960 13637
rect 63632 13588 63674 13628
rect 63714 13588 63756 13628
rect 63796 13588 63838 13628
rect 63878 13588 63920 13628
rect 63592 13579 63960 13588
rect 78712 13628 79080 13637
rect 78752 13588 78794 13628
rect 78834 13588 78876 13628
rect 78916 13588 78958 13628
rect 78998 13588 79040 13628
rect 78712 13579 79080 13588
rect 93832 13628 94200 13637
rect 93872 13588 93914 13628
rect 93954 13588 93996 13628
rect 94036 13588 94078 13628
rect 94118 13588 94160 13628
rect 93832 13579 94200 13588
rect 49712 12872 50080 12881
rect 49752 12832 49794 12872
rect 49834 12832 49876 12872
rect 49916 12832 49958 12872
rect 49998 12832 50040 12872
rect 49712 12823 50080 12832
rect 64832 12872 65200 12881
rect 64872 12832 64914 12872
rect 64954 12832 64996 12872
rect 65036 12832 65078 12872
rect 65118 12832 65160 12872
rect 64832 12823 65200 12832
rect 79952 12872 80320 12881
rect 79992 12832 80034 12872
rect 80074 12832 80116 12872
rect 80156 12832 80198 12872
rect 80238 12832 80280 12872
rect 79952 12823 80320 12832
rect 95072 12872 95440 12881
rect 95112 12832 95154 12872
rect 95194 12832 95236 12872
rect 95276 12832 95318 12872
rect 95358 12832 95400 12872
rect 95072 12823 95440 12832
rect 48472 12116 48840 12125
rect 48512 12076 48554 12116
rect 48594 12076 48636 12116
rect 48676 12076 48718 12116
rect 48758 12076 48800 12116
rect 48472 12067 48840 12076
rect 63592 12116 63960 12125
rect 63632 12076 63674 12116
rect 63714 12076 63756 12116
rect 63796 12076 63838 12116
rect 63878 12076 63920 12116
rect 63592 12067 63960 12076
rect 78712 12116 79080 12125
rect 78752 12076 78794 12116
rect 78834 12076 78876 12116
rect 78916 12076 78958 12116
rect 78998 12076 79040 12116
rect 78712 12067 79080 12076
rect 93832 12116 94200 12125
rect 93872 12076 93914 12116
rect 93954 12076 93996 12116
rect 94036 12076 94078 12116
rect 94118 12076 94160 12116
rect 93832 12067 94200 12076
rect 49712 11360 50080 11369
rect 49752 11320 49794 11360
rect 49834 11320 49876 11360
rect 49916 11320 49958 11360
rect 49998 11320 50040 11360
rect 49712 11311 50080 11320
rect 64832 11360 65200 11369
rect 64872 11320 64914 11360
rect 64954 11320 64996 11360
rect 65036 11320 65078 11360
rect 65118 11320 65160 11360
rect 64832 11311 65200 11320
rect 79952 11360 80320 11369
rect 79992 11320 80034 11360
rect 80074 11320 80116 11360
rect 80156 11320 80198 11360
rect 80238 11320 80280 11360
rect 79952 11311 80320 11320
rect 95072 11360 95440 11369
rect 95112 11320 95154 11360
rect 95194 11320 95236 11360
rect 95276 11320 95318 11360
rect 95358 11320 95400 11360
rect 95072 11311 95440 11320
rect 48472 10604 48840 10613
rect 48512 10564 48554 10604
rect 48594 10564 48636 10604
rect 48676 10564 48718 10604
rect 48758 10564 48800 10604
rect 48472 10555 48840 10564
rect 63592 10604 63960 10613
rect 63632 10564 63674 10604
rect 63714 10564 63756 10604
rect 63796 10564 63838 10604
rect 63878 10564 63920 10604
rect 63592 10555 63960 10564
rect 78712 10604 79080 10613
rect 78752 10564 78794 10604
rect 78834 10564 78876 10604
rect 78916 10564 78958 10604
rect 78998 10564 79040 10604
rect 78712 10555 79080 10564
rect 93832 10604 94200 10613
rect 93872 10564 93914 10604
rect 93954 10564 93996 10604
rect 94036 10564 94078 10604
rect 94118 10564 94160 10604
rect 93832 10555 94200 10564
rect 36747 10268 36789 10277
rect 36747 10228 36748 10268
rect 36788 10228 36789 10268
rect 36747 10219 36789 10228
rect 34592 9848 34960 9857
rect 34632 9808 34674 9848
rect 34714 9808 34756 9848
rect 34796 9808 34838 9848
rect 34878 9808 34920 9848
rect 34592 9799 34960 9808
rect 49712 9848 50080 9857
rect 49752 9808 49794 9848
rect 49834 9808 49876 9848
rect 49916 9808 49958 9848
rect 49998 9808 50040 9848
rect 49712 9799 50080 9808
rect 64832 9848 65200 9857
rect 64872 9808 64914 9848
rect 64954 9808 64996 9848
rect 65036 9808 65078 9848
rect 65118 9808 65160 9848
rect 64832 9799 65200 9808
rect 79952 9848 80320 9857
rect 79992 9808 80034 9848
rect 80074 9808 80116 9848
rect 80156 9808 80198 9848
rect 80238 9808 80280 9848
rect 79952 9799 80320 9808
rect 95072 9848 95440 9857
rect 95112 9808 95154 9848
rect 95194 9808 95236 9848
rect 95276 9808 95318 9848
rect 95358 9808 95400 9848
rect 95072 9799 95440 9808
rect 48472 9092 48840 9101
rect 48512 9052 48554 9092
rect 48594 9052 48636 9092
rect 48676 9052 48718 9092
rect 48758 9052 48800 9092
rect 48472 9043 48840 9052
rect 63592 9092 63960 9101
rect 63632 9052 63674 9092
rect 63714 9052 63756 9092
rect 63796 9052 63838 9092
rect 63878 9052 63920 9092
rect 63592 9043 63960 9052
rect 78712 9092 79080 9101
rect 78752 9052 78794 9092
rect 78834 9052 78876 9092
rect 78916 9052 78958 9092
rect 78998 9052 79040 9092
rect 78712 9043 79080 9052
rect 93832 9092 94200 9101
rect 93872 9052 93914 9092
rect 93954 9052 93996 9092
rect 94036 9052 94078 9092
rect 94118 9052 94160 9092
rect 93832 9043 94200 9052
rect 34592 8336 34960 8345
rect 34632 8296 34674 8336
rect 34714 8296 34756 8336
rect 34796 8296 34838 8336
rect 34878 8296 34920 8336
rect 34592 8287 34960 8296
rect 49712 8336 50080 8345
rect 49752 8296 49794 8336
rect 49834 8296 49876 8336
rect 49916 8296 49958 8336
rect 49998 8296 50040 8336
rect 49712 8287 50080 8296
rect 64832 8336 65200 8345
rect 64872 8296 64914 8336
rect 64954 8296 64996 8336
rect 65036 8296 65078 8336
rect 65118 8296 65160 8336
rect 64832 8287 65200 8296
rect 79952 8336 80320 8345
rect 79992 8296 80034 8336
rect 80074 8296 80116 8336
rect 80156 8296 80198 8336
rect 80238 8296 80280 8336
rect 79952 8287 80320 8296
rect 95072 8336 95440 8345
rect 95112 8296 95154 8336
rect 95194 8296 95236 8336
rect 95276 8296 95318 8336
rect 95358 8296 95400 8336
rect 95072 8287 95440 8296
rect 48472 7580 48840 7589
rect 48512 7540 48554 7580
rect 48594 7540 48636 7580
rect 48676 7540 48718 7580
rect 48758 7540 48800 7580
rect 48472 7531 48840 7540
rect 63592 7580 63960 7589
rect 63632 7540 63674 7580
rect 63714 7540 63756 7580
rect 63796 7540 63838 7580
rect 63878 7540 63920 7580
rect 63592 7531 63960 7540
rect 78712 7580 79080 7589
rect 78752 7540 78794 7580
rect 78834 7540 78876 7580
rect 78916 7540 78958 7580
rect 78998 7540 79040 7580
rect 78712 7531 79080 7540
rect 93832 7580 94200 7589
rect 93872 7540 93914 7580
rect 93954 7540 93996 7580
rect 94036 7540 94078 7580
rect 94118 7540 94160 7580
rect 93832 7531 94200 7540
rect 34592 6824 34960 6833
rect 34632 6784 34674 6824
rect 34714 6784 34756 6824
rect 34796 6784 34838 6824
rect 34878 6784 34920 6824
rect 34592 6775 34960 6784
rect 49712 6824 50080 6833
rect 49752 6784 49794 6824
rect 49834 6784 49876 6824
rect 49916 6784 49958 6824
rect 49998 6784 50040 6824
rect 49712 6775 50080 6784
rect 64832 6824 65200 6833
rect 64872 6784 64914 6824
rect 64954 6784 64996 6824
rect 65036 6784 65078 6824
rect 65118 6784 65160 6824
rect 64832 6775 65200 6784
rect 79952 6824 80320 6833
rect 79992 6784 80034 6824
rect 80074 6784 80116 6824
rect 80156 6784 80198 6824
rect 80238 6784 80280 6824
rect 79952 6775 80320 6784
rect 95072 6824 95440 6833
rect 95112 6784 95154 6824
rect 95194 6784 95236 6824
rect 95276 6784 95318 6824
rect 95358 6784 95400 6824
rect 95072 6775 95440 6784
rect 48472 6068 48840 6077
rect 48512 6028 48554 6068
rect 48594 6028 48636 6068
rect 48676 6028 48718 6068
rect 48758 6028 48800 6068
rect 48472 6019 48840 6028
rect 63592 6068 63960 6077
rect 63632 6028 63674 6068
rect 63714 6028 63756 6068
rect 63796 6028 63838 6068
rect 63878 6028 63920 6068
rect 63592 6019 63960 6028
rect 78712 6068 79080 6077
rect 78752 6028 78794 6068
rect 78834 6028 78876 6068
rect 78916 6028 78958 6068
rect 78998 6028 79040 6068
rect 78712 6019 79080 6028
rect 93832 6068 94200 6077
rect 93872 6028 93914 6068
rect 93954 6028 93996 6068
rect 94036 6028 94078 6068
rect 94118 6028 94160 6068
rect 93832 6019 94200 6028
rect 34592 5312 34960 5321
rect 34632 5272 34674 5312
rect 34714 5272 34756 5312
rect 34796 5272 34838 5312
rect 34878 5272 34920 5312
rect 34592 5263 34960 5272
rect 49712 5312 50080 5321
rect 49752 5272 49794 5312
rect 49834 5272 49876 5312
rect 49916 5272 49958 5312
rect 49998 5272 50040 5312
rect 49712 5263 50080 5272
rect 64832 5312 65200 5321
rect 64872 5272 64914 5312
rect 64954 5272 64996 5312
rect 65036 5272 65078 5312
rect 65118 5272 65160 5312
rect 64832 5263 65200 5272
rect 79952 5312 80320 5321
rect 79992 5272 80034 5312
rect 80074 5272 80116 5312
rect 80156 5272 80198 5312
rect 80238 5272 80280 5312
rect 79952 5263 80320 5272
rect 95072 5312 95440 5321
rect 95112 5272 95154 5312
rect 95194 5272 95236 5312
rect 95276 5272 95318 5312
rect 95358 5272 95400 5312
rect 95072 5263 95440 5272
rect 48472 4556 48840 4565
rect 48512 4516 48554 4556
rect 48594 4516 48636 4556
rect 48676 4516 48718 4556
rect 48758 4516 48800 4556
rect 48472 4507 48840 4516
rect 63592 4556 63960 4565
rect 63632 4516 63674 4556
rect 63714 4516 63756 4556
rect 63796 4516 63838 4556
rect 63878 4516 63920 4556
rect 63592 4507 63960 4516
rect 78712 4556 79080 4565
rect 78752 4516 78794 4556
rect 78834 4516 78876 4556
rect 78916 4516 78958 4556
rect 78998 4516 79040 4556
rect 78712 4507 79080 4516
rect 93832 4556 94200 4565
rect 93872 4516 93914 4556
rect 93954 4516 93996 4556
rect 94036 4516 94078 4556
rect 94118 4516 94160 4556
rect 93832 4507 94200 4516
rect 34443 4220 34485 4229
rect 34443 4180 34444 4220
rect 34484 4180 34485 4220
rect 34443 4171 34485 4180
rect 4352 3800 4720 3809
rect 4392 3760 4434 3800
rect 4474 3760 4516 3800
rect 4556 3760 4598 3800
rect 4638 3760 4680 3800
rect 4352 3751 4720 3760
rect 19472 3800 19840 3809
rect 19512 3760 19554 3800
rect 19594 3760 19636 3800
rect 19676 3760 19718 3800
rect 19758 3760 19800 3800
rect 19472 3751 19840 3760
rect 34592 3800 34960 3809
rect 34632 3760 34674 3800
rect 34714 3760 34756 3800
rect 34796 3760 34838 3800
rect 34878 3760 34920 3800
rect 34592 3751 34960 3760
rect 49712 3800 50080 3809
rect 49752 3760 49794 3800
rect 49834 3760 49876 3800
rect 49916 3760 49958 3800
rect 49998 3760 50040 3800
rect 49712 3751 50080 3760
rect 64832 3800 65200 3809
rect 64872 3760 64914 3800
rect 64954 3760 64996 3800
rect 65036 3760 65078 3800
rect 65118 3760 65160 3800
rect 64832 3751 65200 3760
rect 79952 3800 80320 3809
rect 79992 3760 80034 3800
rect 80074 3760 80116 3800
rect 80156 3760 80198 3800
rect 80238 3760 80280 3800
rect 79952 3751 80320 3760
rect 95072 3800 95440 3809
rect 95112 3760 95154 3800
rect 95194 3760 95236 3800
rect 95276 3760 95318 3800
rect 95358 3760 95400 3800
rect 95072 3751 95440 3760
rect 884 3340 1172 3380
rect 844 3331 884 3340
rect 3112 3044 3480 3053
rect 3152 3004 3194 3044
rect 3234 3004 3276 3044
rect 3316 3004 3358 3044
rect 3398 3004 3440 3044
rect 3112 2995 3480 3004
rect 18232 3044 18600 3053
rect 18272 3004 18314 3044
rect 18354 3004 18396 3044
rect 18436 3004 18478 3044
rect 18518 3004 18560 3044
rect 18232 2995 18600 3004
rect 33352 3044 33720 3053
rect 33392 3004 33434 3044
rect 33474 3004 33516 3044
rect 33556 3004 33598 3044
rect 33638 3004 33680 3044
rect 33352 2995 33720 3004
rect 48472 3044 48840 3053
rect 48512 3004 48554 3044
rect 48594 3004 48636 3044
rect 48676 3004 48718 3044
rect 48758 3004 48800 3044
rect 48472 2995 48840 3004
rect 63592 3044 63960 3053
rect 63632 3004 63674 3044
rect 63714 3004 63756 3044
rect 63796 3004 63838 3044
rect 63878 3004 63920 3044
rect 63592 2995 63960 3004
rect 78712 3044 79080 3053
rect 78752 3004 78794 3044
rect 78834 3004 78876 3044
rect 78916 3004 78958 3044
rect 78998 3004 79040 3044
rect 78712 2995 79080 3004
rect 93832 3044 94200 3053
rect 93872 3004 93914 3044
rect 93954 3004 93996 3044
rect 94036 3004 94078 3044
rect 94118 3004 94160 3044
rect 93832 2995 94200 3004
rect 844 2708 884 2717
rect 748 2668 844 2708
rect 844 2659 884 2668
rect 652 2456 692 2465
rect 652 2297 692 2416
rect 651 2288 693 2297
rect 651 2248 652 2288
rect 692 2248 693 2288
rect 651 2239 693 2248
rect 4352 2288 4720 2297
rect 4392 2248 4434 2288
rect 4474 2248 4516 2288
rect 4556 2248 4598 2288
rect 4638 2248 4680 2288
rect 4352 2239 4720 2248
rect 19472 2288 19840 2297
rect 19512 2248 19554 2288
rect 19594 2248 19636 2288
rect 19676 2248 19718 2288
rect 19758 2248 19800 2288
rect 19472 2239 19840 2248
rect 34592 2288 34960 2297
rect 34632 2248 34674 2288
rect 34714 2248 34756 2288
rect 34796 2248 34838 2288
rect 34878 2248 34920 2288
rect 34592 2239 34960 2248
rect 49712 2288 50080 2297
rect 49752 2248 49794 2288
rect 49834 2248 49876 2288
rect 49916 2248 49958 2288
rect 49998 2248 50040 2288
rect 49712 2239 50080 2248
rect 64832 2288 65200 2297
rect 64872 2248 64914 2288
rect 64954 2248 64996 2288
rect 65036 2248 65078 2288
rect 65118 2248 65160 2288
rect 64832 2239 65200 2248
rect 79952 2288 80320 2297
rect 79992 2248 80034 2288
rect 80074 2248 80116 2288
rect 80156 2248 80198 2288
rect 80238 2248 80280 2288
rect 79952 2239 80320 2248
rect 95072 2288 95440 2297
rect 95112 2248 95154 2288
rect 95194 2248 95236 2288
rect 95276 2248 95318 2288
rect 95358 2248 95400 2288
rect 95072 2239 95440 2248
rect 3112 1532 3480 1541
rect 3152 1492 3194 1532
rect 3234 1492 3276 1532
rect 3316 1492 3358 1532
rect 3398 1492 3440 1532
rect 3112 1483 3480 1492
rect 18232 1532 18600 1541
rect 18272 1492 18314 1532
rect 18354 1492 18396 1532
rect 18436 1492 18478 1532
rect 18518 1492 18560 1532
rect 18232 1483 18600 1492
rect 33352 1532 33720 1541
rect 33392 1492 33434 1532
rect 33474 1492 33516 1532
rect 33556 1492 33598 1532
rect 33638 1492 33680 1532
rect 33352 1483 33720 1492
rect 48472 1532 48840 1541
rect 48512 1492 48554 1532
rect 48594 1492 48636 1532
rect 48676 1492 48718 1532
rect 48758 1492 48800 1532
rect 48472 1483 48840 1492
rect 63592 1532 63960 1541
rect 63632 1492 63674 1532
rect 63714 1492 63756 1532
rect 63796 1492 63838 1532
rect 63878 1492 63920 1532
rect 63592 1483 63960 1492
rect 78712 1532 79080 1541
rect 78752 1492 78794 1532
rect 78834 1492 78876 1532
rect 78916 1492 78958 1532
rect 78998 1492 79040 1532
rect 78712 1483 79080 1492
rect 93832 1532 94200 1541
rect 93872 1492 93914 1532
rect 93954 1492 93996 1532
rect 94036 1492 94078 1532
rect 94118 1492 94160 1532
rect 93832 1483 94200 1492
rect 4352 776 4720 785
rect 4392 736 4434 776
rect 4474 736 4516 776
rect 4556 736 4598 776
rect 4638 736 4680 776
rect 4352 727 4720 736
rect 19472 776 19840 785
rect 19512 736 19554 776
rect 19594 736 19636 776
rect 19676 736 19718 776
rect 19758 736 19800 776
rect 19472 727 19840 736
rect 34592 776 34960 785
rect 34632 736 34674 776
rect 34714 736 34756 776
rect 34796 736 34838 776
rect 34878 736 34920 776
rect 34592 727 34960 736
rect 49712 776 50080 785
rect 49752 736 49794 776
rect 49834 736 49876 776
rect 49916 736 49958 776
rect 49998 736 50040 776
rect 49712 727 50080 736
rect 64832 776 65200 785
rect 64872 736 64914 776
rect 64954 736 64996 776
rect 65036 736 65078 776
rect 65118 736 65160 776
rect 64832 727 65200 736
rect 79952 776 80320 785
rect 79992 736 80034 776
rect 80074 736 80116 776
rect 80156 736 80198 776
rect 80238 736 80280 776
rect 79952 727 80320 736
rect 95072 776 95440 785
rect 95112 736 95154 776
rect 95194 736 95236 776
rect 95276 736 95318 776
rect 95358 736 95400 776
rect 95072 727 95440 736
<< via2 >>
rect 4352 38536 4392 38576
rect 4434 38536 4474 38576
rect 4516 38536 4556 38576
rect 4598 38536 4638 38576
rect 4680 38536 4720 38576
rect 19472 38536 19512 38576
rect 19554 38536 19594 38576
rect 19636 38536 19676 38576
rect 19718 38536 19758 38576
rect 19800 38536 19840 38576
rect 34592 38536 34632 38576
rect 34674 38536 34714 38576
rect 34756 38536 34796 38576
rect 34838 38536 34878 38576
rect 34920 38536 34960 38576
rect 49712 38536 49752 38576
rect 49794 38536 49834 38576
rect 49876 38536 49916 38576
rect 49958 38536 49998 38576
rect 50040 38536 50080 38576
rect 64832 38536 64872 38576
rect 64914 38536 64954 38576
rect 64996 38536 65036 38576
rect 65078 38536 65118 38576
rect 65160 38536 65200 38576
rect 79952 38536 79992 38576
rect 80034 38536 80074 38576
rect 80116 38536 80156 38576
rect 80198 38536 80238 38576
rect 80280 38536 80320 38576
rect 95072 38536 95112 38576
rect 95154 38536 95194 38576
rect 95236 38536 95276 38576
rect 95318 38536 95358 38576
rect 95400 38536 95440 38576
rect 3112 37780 3152 37820
rect 3194 37780 3234 37820
rect 3276 37780 3316 37820
rect 3358 37780 3398 37820
rect 3440 37780 3480 37820
rect 18232 37780 18272 37820
rect 18314 37780 18354 37820
rect 18396 37780 18436 37820
rect 18478 37780 18518 37820
rect 18560 37780 18600 37820
rect 33352 37780 33392 37820
rect 33434 37780 33474 37820
rect 33516 37780 33556 37820
rect 33598 37780 33638 37820
rect 33680 37780 33720 37820
rect 48472 37780 48512 37820
rect 48554 37780 48594 37820
rect 48636 37780 48676 37820
rect 48718 37780 48758 37820
rect 48800 37780 48840 37820
rect 63592 37780 63632 37820
rect 63674 37780 63714 37820
rect 63756 37780 63796 37820
rect 63838 37780 63878 37820
rect 63920 37780 63960 37820
rect 78712 37780 78752 37820
rect 78794 37780 78834 37820
rect 78876 37780 78916 37820
rect 78958 37780 78998 37820
rect 79040 37780 79080 37820
rect 93832 37780 93872 37820
rect 93914 37780 93954 37820
rect 93996 37780 94036 37820
rect 94078 37780 94118 37820
rect 94160 37780 94200 37820
rect 268 37528 308 37568
rect 76 36688 116 36728
rect 4352 37024 4392 37064
rect 4434 37024 4474 37064
rect 4516 37024 4556 37064
rect 4598 37024 4638 37064
rect 4680 37024 4720 37064
rect 19472 37024 19512 37064
rect 19554 37024 19594 37064
rect 19636 37024 19676 37064
rect 19718 37024 19758 37064
rect 19800 37024 19840 37064
rect 34592 37024 34632 37064
rect 34674 37024 34714 37064
rect 34756 37024 34796 37064
rect 34838 37024 34878 37064
rect 34920 37024 34960 37064
rect 49712 37024 49752 37064
rect 49794 37024 49834 37064
rect 49876 37024 49916 37064
rect 49958 37024 49998 37064
rect 50040 37024 50080 37064
rect 64832 37024 64872 37064
rect 64914 37024 64954 37064
rect 64996 37024 65036 37064
rect 65078 37024 65118 37064
rect 65160 37024 65200 37064
rect 79952 37024 79992 37064
rect 80034 37024 80074 37064
rect 80116 37024 80156 37064
rect 80198 37024 80238 37064
rect 80280 37024 80320 37064
rect 95072 37024 95112 37064
rect 95154 37024 95194 37064
rect 95236 37024 95276 37064
rect 95318 37024 95358 37064
rect 95400 37024 95440 37064
rect 3112 36268 3152 36308
rect 3194 36268 3234 36308
rect 3276 36268 3316 36308
rect 3358 36268 3398 36308
rect 3440 36268 3480 36308
rect 18232 36268 18272 36308
rect 18314 36268 18354 36308
rect 18396 36268 18436 36308
rect 18478 36268 18518 36308
rect 18560 36268 18600 36308
rect 33352 36268 33392 36308
rect 33434 36268 33474 36308
rect 33516 36268 33556 36308
rect 33598 36268 33638 36308
rect 33680 36268 33720 36308
rect 48472 36268 48512 36308
rect 48554 36268 48594 36308
rect 48636 36268 48676 36308
rect 48718 36268 48758 36308
rect 48800 36268 48840 36308
rect 63592 36268 63632 36308
rect 63674 36268 63714 36308
rect 63756 36268 63796 36308
rect 63838 36268 63878 36308
rect 63920 36268 63960 36308
rect 78712 36268 78752 36308
rect 78794 36268 78834 36308
rect 78876 36268 78916 36308
rect 78958 36268 78998 36308
rect 79040 36268 79080 36308
rect 93832 36268 93872 36308
rect 93914 36268 93954 36308
rect 93996 36268 94036 36308
rect 94078 36268 94118 36308
rect 94160 36268 94200 36308
rect 4352 35512 4392 35552
rect 4434 35512 4474 35552
rect 4516 35512 4556 35552
rect 4598 35512 4638 35552
rect 4680 35512 4720 35552
rect 19472 35512 19512 35552
rect 19554 35512 19594 35552
rect 19636 35512 19676 35552
rect 19718 35512 19758 35552
rect 19800 35512 19840 35552
rect 34592 35512 34632 35552
rect 34674 35512 34714 35552
rect 34756 35512 34796 35552
rect 34838 35512 34878 35552
rect 34920 35512 34960 35552
rect 49712 35512 49752 35552
rect 49794 35512 49834 35552
rect 49876 35512 49916 35552
rect 49958 35512 49998 35552
rect 50040 35512 50080 35552
rect 64832 35512 64872 35552
rect 64914 35512 64954 35552
rect 64996 35512 65036 35552
rect 65078 35512 65118 35552
rect 65160 35512 65200 35552
rect 79952 35512 79992 35552
rect 80034 35512 80074 35552
rect 80116 35512 80156 35552
rect 80198 35512 80238 35552
rect 80280 35512 80320 35552
rect 95072 35512 95112 35552
rect 95154 35512 95194 35552
rect 95236 35512 95276 35552
rect 95318 35512 95358 35552
rect 95400 35512 95440 35552
rect 844 35176 884 35216
rect 23500 35176 23540 35216
rect 652 35008 692 35048
rect 3112 34756 3152 34796
rect 3194 34756 3234 34796
rect 3276 34756 3316 34796
rect 3358 34756 3398 34796
rect 3440 34756 3480 34796
rect 18232 34756 18272 34796
rect 18314 34756 18354 34796
rect 18396 34756 18436 34796
rect 18478 34756 18518 34796
rect 18560 34756 18600 34796
rect 844 34336 884 34376
rect 652 34168 692 34208
rect 4352 34000 4392 34040
rect 4434 34000 4474 34040
rect 4516 34000 4556 34040
rect 4598 34000 4638 34040
rect 4680 34000 4720 34040
rect 19472 34000 19512 34040
rect 19554 34000 19594 34040
rect 19636 34000 19676 34040
rect 19718 34000 19758 34040
rect 19800 34000 19840 34040
rect 844 33664 884 33704
rect 652 33328 692 33368
rect 3112 33244 3152 33284
rect 3194 33244 3234 33284
rect 3276 33244 3316 33284
rect 3358 33244 3398 33284
rect 3440 33244 3480 33284
rect 18232 33244 18272 33284
rect 18314 33244 18354 33284
rect 18396 33244 18436 33284
rect 18478 33244 18518 33284
rect 18560 33244 18600 33284
rect 844 32824 884 32864
rect 652 32488 692 32528
rect 4352 32488 4392 32528
rect 4434 32488 4474 32528
rect 4516 32488 4556 32528
rect 4598 32488 4638 32528
rect 4680 32488 4720 32528
rect 19472 32488 19512 32528
rect 19554 32488 19594 32528
rect 19636 32488 19676 32528
rect 19718 32488 19758 32528
rect 19800 32488 19840 32528
rect 652 31648 692 31688
rect 652 30808 692 30848
rect 652 30052 692 30092
rect 652 29128 692 29168
rect 652 28288 692 28328
rect 844 28288 884 28328
rect 748 27784 788 27824
rect 652 27448 692 27488
rect 940 27448 980 27488
rect 3112 31732 3152 31772
rect 3194 31732 3234 31772
rect 3276 31732 3316 31772
rect 3358 31732 3398 31772
rect 3440 31732 3480 31772
rect 18232 31732 18272 31772
rect 18314 31732 18354 31772
rect 18396 31732 18436 31772
rect 18478 31732 18518 31772
rect 18560 31732 18600 31772
rect 22636 31312 22676 31352
rect 4352 30976 4392 31016
rect 4434 30976 4474 31016
rect 4516 30976 4556 31016
rect 4598 30976 4638 31016
rect 4680 30976 4720 31016
rect 19472 30976 19512 31016
rect 19554 30976 19594 31016
rect 19636 30976 19676 31016
rect 19718 30976 19758 31016
rect 19800 30976 19840 31016
rect 3112 30220 3152 30260
rect 3194 30220 3234 30260
rect 3276 30220 3316 30260
rect 3358 30220 3398 30260
rect 3440 30220 3480 30260
rect 18232 30220 18272 30260
rect 18314 30220 18354 30260
rect 18396 30220 18436 30260
rect 18478 30220 18518 30260
rect 18560 30220 18600 30260
rect 1132 29800 1172 29840
rect 19948 29800 19988 29840
rect 4352 29464 4392 29504
rect 4434 29464 4474 29504
rect 4516 29464 4556 29504
rect 4598 29464 4638 29504
rect 4680 29464 4720 29504
rect 19472 29464 19512 29504
rect 19554 29464 19594 29504
rect 19636 29464 19676 29504
rect 19718 29464 19758 29504
rect 19800 29464 19840 29504
rect 3112 28708 3152 28748
rect 3194 28708 3234 28748
rect 3276 28708 3316 28748
rect 3358 28708 3398 28748
rect 3440 28708 3480 28748
rect 15340 28288 15380 28328
rect 4352 27952 4392 27992
rect 4434 27952 4474 27992
rect 4516 27952 4556 27992
rect 4598 27952 4638 27992
rect 4680 27952 4720 27992
rect 3112 27196 3152 27236
rect 3194 27196 3234 27236
rect 3276 27196 3316 27236
rect 3358 27196 3398 27236
rect 3440 27196 3480 27236
rect 652 26608 692 26648
rect 268 26188 308 26228
rect 172 21568 212 21608
rect 652 25768 692 25808
rect 652 24928 692 24968
rect 652 24088 692 24128
rect 652 23248 692 23288
rect 652 21652 692 21692
rect 652 20728 692 20768
rect 1036 26944 1076 26984
rect 14860 26608 14900 26648
rect 4352 26440 4392 26480
rect 4434 26440 4474 26480
rect 4516 26440 4556 26480
rect 4598 26440 4638 26480
rect 4680 26440 4720 26480
rect 18232 28708 18272 28748
rect 18314 28708 18354 28748
rect 18396 28708 18436 28748
rect 18478 28708 18518 28748
rect 18560 28708 18600 28748
rect 18220 28036 18260 28076
rect 17260 27616 17300 27656
rect 18124 27616 18164 27656
rect 16108 26356 16148 26396
rect 16588 26356 16628 26396
rect 19472 27952 19512 27992
rect 19554 27952 19594 27992
rect 19636 27952 19676 27992
rect 19718 27952 19758 27992
rect 19800 27952 19840 27992
rect 21772 31228 21812 31268
rect 21388 28540 21428 28580
rect 20044 27784 20084 27824
rect 18508 27616 18548 27656
rect 18232 27196 18272 27236
rect 18314 27196 18354 27236
rect 18396 27196 18436 27236
rect 18478 27196 18518 27236
rect 18560 27196 18600 27236
rect 3112 25684 3152 25724
rect 3194 25684 3234 25724
rect 3276 25684 3316 25724
rect 3358 25684 3398 25724
rect 3440 25684 3480 25724
rect 940 25432 980 25472
rect 844 23752 884 23792
rect 940 20728 980 20768
rect 748 19972 788 20012
rect 652 19888 692 19928
rect 556 19804 596 19844
rect 4352 24928 4392 24968
rect 4434 24928 4474 24968
rect 4516 24928 4556 24968
rect 4598 24928 4638 24968
rect 4680 24928 4720 24968
rect 3112 24172 3152 24212
rect 3194 24172 3234 24212
rect 3276 24172 3316 24212
rect 3358 24172 3398 24212
rect 3440 24172 3480 24212
rect 4352 23416 4392 23456
rect 4434 23416 4474 23456
rect 4516 23416 4556 23456
rect 4598 23416 4638 23456
rect 4680 23416 4720 23456
rect 18232 25684 18272 25724
rect 18314 25684 18354 25724
rect 18396 25684 18436 25724
rect 18478 25684 18518 25724
rect 18560 25684 18600 25724
rect 18232 24172 18272 24212
rect 18314 24172 18354 24212
rect 18396 24172 18436 24212
rect 18478 24172 18518 24212
rect 18560 24172 18600 24212
rect 21484 27784 21524 27824
rect 20236 27616 20276 27656
rect 20140 27448 20180 27488
rect 19948 26944 19988 26984
rect 20236 26860 20276 26900
rect 20428 26860 20468 26900
rect 20140 26776 20180 26816
rect 20620 26776 20660 26816
rect 20332 26608 20372 26648
rect 19472 26440 19512 26480
rect 19554 26440 19594 26480
rect 19636 26440 19676 26480
rect 19718 26440 19758 26480
rect 19800 26440 19840 26480
rect 21580 27700 21620 27740
rect 21676 27448 21716 27488
rect 21772 26776 21812 26816
rect 19472 24928 19512 24968
rect 19554 24928 19594 24968
rect 19636 24928 19676 24968
rect 19718 24928 19758 24968
rect 19800 24928 19840 24968
rect 15244 23080 15284 23120
rect 3112 22660 3152 22700
rect 3194 22660 3234 22700
rect 3276 22660 3316 22700
rect 3358 22660 3398 22700
rect 3440 22660 3480 22700
rect 4352 21904 4392 21944
rect 4434 21904 4474 21944
rect 4516 21904 4556 21944
rect 4598 21904 4638 21944
rect 4680 21904 4720 21944
rect 3112 21148 3152 21188
rect 3194 21148 3234 21188
rect 3276 21148 3316 21188
rect 3358 21148 3398 21188
rect 3440 21148 3480 21188
rect 1132 20476 1172 20516
rect 1036 19468 1076 19508
rect 652 19048 692 19088
rect 652 18208 692 18248
rect 652 17368 692 17408
rect 652 16528 692 16568
rect 556 15688 596 15728
rect 940 15268 980 15308
rect 652 14848 692 14888
rect 652 14008 692 14048
rect 652 13168 692 13208
rect 844 13000 884 13040
rect 652 12328 692 12368
rect 748 12160 788 12200
rect 652 11488 692 11528
rect 652 10732 692 10772
rect 652 9808 692 9848
rect 652 8968 692 9008
rect 844 10900 884 10940
rect 844 10228 884 10268
rect 844 9388 884 9428
rect 1036 11992 1076 12032
rect 652 8128 692 8168
rect 652 7288 692 7328
rect 652 6448 692 6488
rect 652 5608 692 5648
rect 652 4768 692 4808
rect 652 3928 692 3968
rect 652 3172 692 3212
rect 844 7204 884 7244
rect 844 5692 884 5732
rect 844 4852 884 4892
rect 844 4180 884 4220
rect 4352 20392 4392 20432
rect 4434 20392 4474 20432
rect 4516 20392 4556 20432
rect 4598 20392 4638 20432
rect 4680 20392 4720 20432
rect 17356 22072 17396 22112
rect 17740 20728 17780 20768
rect 14956 20140 14996 20180
rect 15436 20140 15476 20180
rect 15916 19972 15956 20012
rect 15628 19888 15668 19928
rect 3112 19636 3152 19676
rect 3194 19636 3234 19676
rect 3276 19636 3316 19676
rect 3358 19636 3398 19676
rect 3440 19636 3480 19676
rect 15916 19216 15956 19256
rect 16108 19216 16148 19256
rect 15724 19132 15764 19172
rect 4352 18880 4392 18920
rect 4434 18880 4474 18920
rect 4516 18880 4556 18920
rect 4598 18880 4638 18920
rect 4680 18880 4720 18920
rect 3112 18124 3152 18164
rect 3194 18124 3234 18164
rect 3276 18124 3316 18164
rect 3358 18124 3398 18164
rect 3440 18124 3480 18164
rect 4352 17368 4392 17408
rect 4434 17368 4474 17408
rect 4516 17368 4556 17408
rect 4598 17368 4638 17408
rect 4680 17368 4720 17408
rect 18028 19468 18068 19508
rect 16204 17704 16244 17744
rect 17644 17704 17684 17744
rect 3112 16612 3152 16652
rect 3194 16612 3234 16652
rect 3276 16612 3316 16652
rect 3358 16612 3398 16652
rect 3440 16612 3480 16652
rect 4352 15856 4392 15896
rect 4434 15856 4474 15896
rect 4516 15856 4556 15896
rect 4598 15856 4638 15896
rect 4680 15856 4720 15896
rect 3112 15100 3152 15140
rect 3194 15100 3234 15140
rect 3276 15100 3316 15140
rect 3358 15100 3398 15140
rect 3440 15100 3480 15140
rect 4352 14344 4392 14384
rect 4434 14344 4474 14384
rect 4516 14344 4556 14384
rect 4598 14344 4638 14384
rect 4680 14344 4720 14384
rect 3112 13588 3152 13628
rect 3194 13588 3234 13628
rect 3276 13588 3316 13628
rect 3358 13588 3398 13628
rect 3440 13588 3480 13628
rect 4352 12832 4392 12872
rect 4434 12832 4474 12872
rect 4516 12832 4556 12872
rect 4598 12832 4638 12872
rect 4680 12832 4720 12872
rect 16684 15520 16724 15560
rect 17836 15688 17876 15728
rect 19472 23416 19512 23456
rect 19554 23416 19594 23456
rect 19636 23416 19676 23456
rect 19718 23416 19758 23456
rect 19800 23416 19840 23456
rect 22060 28540 22100 28580
rect 22444 28288 22484 28328
rect 22348 27784 22388 27824
rect 22540 27700 22580 27740
rect 23212 28288 23252 28328
rect 23404 28288 23444 28328
rect 33352 34756 33392 34796
rect 33434 34756 33474 34796
rect 33516 34756 33556 34796
rect 33598 34756 33638 34796
rect 33680 34756 33720 34796
rect 48472 34756 48512 34796
rect 48554 34756 48594 34796
rect 48636 34756 48676 34796
rect 48718 34756 48758 34796
rect 48800 34756 48840 34796
rect 63592 34756 63632 34796
rect 63674 34756 63714 34796
rect 63756 34756 63796 34796
rect 63838 34756 63878 34796
rect 63920 34756 63960 34796
rect 78712 34756 78752 34796
rect 78794 34756 78834 34796
rect 78876 34756 78916 34796
rect 78958 34756 78998 34796
rect 79040 34756 79080 34796
rect 93832 34756 93872 34796
rect 93914 34756 93954 34796
rect 93996 34756 94036 34796
rect 94078 34756 94118 34796
rect 94160 34756 94200 34796
rect 29356 34336 29396 34376
rect 29068 32824 29108 32864
rect 27052 31900 27092 31940
rect 23788 31144 23828 31184
rect 26764 30640 26804 30680
rect 23500 28120 23540 28160
rect 26860 28120 26900 28160
rect 23404 28036 23444 28076
rect 23308 27784 23348 27824
rect 23404 27700 23444 27740
rect 26572 27700 26612 27740
rect 26380 27616 26420 27656
rect 23596 27364 23636 27404
rect 25804 26860 25844 26900
rect 26380 26860 26420 26900
rect 22636 26356 22676 26396
rect 26956 27616 26996 27656
rect 25996 26020 26036 26060
rect 26380 26020 26420 26060
rect 26860 26020 26900 26060
rect 26380 25516 26420 25556
rect 22636 24592 22676 24632
rect 23020 24592 23060 24632
rect 18232 22660 18272 22700
rect 18314 22660 18354 22700
rect 18396 22660 18436 22700
rect 18478 22660 18518 22700
rect 18560 22660 18600 22700
rect 18232 21148 18272 21188
rect 18314 21148 18354 21188
rect 18396 21148 18436 21188
rect 18478 21148 18518 21188
rect 18560 21148 18600 21188
rect 19756 23080 19796 23120
rect 19472 21904 19512 21944
rect 19554 21904 19594 21944
rect 19636 21904 19676 21944
rect 19718 21904 19758 21944
rect 19800 21904 19840 21944
rect 18232 19636 18272 19676
rect 18314 19636 18354 19676
rect 18396 19636 18436 19676
rect 18478 19636 18518 19676
rect 18560 19636 18600 19676
rect 19180 19300 19220 19340
rect 19084 19132 19124 19172
rect 19564 20728 19604 20768
rect 20140 20728 20180 20768
rect 19472 20392 19512 20432
rect 19554 20392 19594 20432
rect 19636 20392 19676 20432
rect 19718 20392 19758 20432
rect 19800 20392 19840 20432
rect 20140 20140 20180 20180
rect 19468 20056 19508 20096
rect 19468 19468 19508 19508
rect 19372 19300 19412 19340
rect 19660 19216 19700 19256
rect 18232 18124 18272 18164
rect 18314 18124 18354 18164
rect 18396 18124 18436 18164
rect 18478 18124 18518 18164
rect 18560 18124 18600 18164
rect 19472 18880 19512 18920
rect 19554 18880 19594 18920
rect 19636 18880 19676 18920
rect 19718 18880 19758 18920
rect 19800 18880 19840 18920
rect 19372 17704 19412 17744
rect 19472 17368 19512 17408
rect 19554 17368 19594 17408
rect 19636 17368 19676 17408
rect 19718 17368 19758 17408
rect 19800 17368 19840 17408
rect 18232 16612 18272 16652
rect 18314 16612 18354 16652
rect 18396 16612 18436 16652
rect 18478 16612 18518 16652
rect 18560 16612 18600 16652
rect 19472 15856 19512 15896
rect 19554 15856 19594 15896
rect 19636 15856 19676 15896
rect 19718 15856 19758 15896
rect 19800 15856 19840 15896
rect 18220 15688 18260 15728
rect 21868 23080 21908 23120
rect 21772 22828 21812 22868
rect 23404 22156 23444 22196
rect 22636 20728 22676 20768
rect 22060 20308 22100 20348
rect 21772 20140 21812 20180
rect 22348 20140 22388 20180
rect 21100 19300 21140 19340
rect 21388 20056 21428 20096
rect 21868 20056 21908 20096
rect 21388 19888 21428 19928
rect 21292 19216 21332 19256
rect 21100 18628 21140 18668
rect 21388 17956 21428 17996
rect 22060 17956 22100 17996
rect 22252 17956 22292 17996
rect 18988 15520 19028 15560
rect 20620 15520 20660 15560
rect 18412 15436 18452 15476
rect 18508 15352 18548 15392
rect 18892 15352 18932 15392
rect 18700 15268 18740 15308
rect 18232 15100 18272 15140
rect 18314 15100 18354 15140
rect 18396 15100 18436 15140
rect 18478 15100 18518 15140
rect 18560 15100 18600 15140
rect 15820 12496 15860 12536
rect 3112 12076 3152 12116
rect 3194 12076 3234 12116
rect 3276 12076 3316 12116
rect 3358 12076 3398 12116
rect 3440 12076 3480 12116
rect 4352 11320 4392 11360
rect 4434 11320 4474 11360
rect 4516 11320 4556 11360
rect 4598 11320 4638 11360
rect 4680 11320 4720 11360
rect 18232 13588 18272 13628
rect 18314 13588 18354 13628
rect 18396 13588 18436 13628
rect 18478 13588 18518 13628
rect 18560 13588 18600 13628
rect 18124 12496 18164 12536
rect 18232 12076 18272 12116
rect 18314 12076 18354 12116
rect 18396 12076 18436 12116
rect 18478 12076 18518 12116
rect 18560 12076 18600 12116
rect 18028 10900 18068 10940
rect 3112 10564 3152 10604
rect 3194 10564 3234 10604
rect 3276 10564 3316 10604
rect 3358 10564 3398 10604
rect 3440 10564 3480 10604
rect 18232 10564 18272 10604
rect 18314 10564 18354 10604
rect 18396 10564 18436 10604
rect 18478 10564 18518 10604
rect 18560 10564 18600 10604
rect 4352 9808 4392 9848
rect 4434 9808 4474 9848
rect 4516 9808 4556 9848
rect 4598 9808 4638 9848
rect 4680 9808 4720 9848
rect 3112 9052 3152 9092
rect 3194 9052 3234 9092
rect 3276 9052 3316 9092
rect 3358 9052 3398 9092
rect 3440 9052 3480 9092
rect 18232 9052 18272 9092
rect 18314 9052 18354 9092
rect 18396 9052 18436 9092
rect 18478 9052 18518 9092
rect 18560 9052 18600 9092
rect 4352 8296 4392 8336
rect 4434 8296 4474 8336
rect 4516 8296 4556 8336
rect 4598 8296 4638 8336
rect 4680 8296 4720 8336
rect 3112 7540 3152 7580
rect 3194 7540 3234 7580
rect 3276 7540 3316 7580
rect 3358 7540 3398 7580
rect 3440 7540 3480 7580
rect 18232 7540 18272 7580
rect 18314 7540 18354 7580
rect 18396 7540 18436 7580
rect 18478 7540 18518 7580
rect 18560 7540 18600 7580
rect 4352 6784 4392 6824
rect 4434 6784 4474 6824
rect 4516 6784 4556 6824
rect 4598 6784 4638 6824
rect 4680 6784 4720 6824
rect 22540 19132 22580 19172
rect 22444 18628 22484 18668
rect 22444 18292 22484 18332
rect 22732 20308 22772 20348
rect 22924 20644 22964 20684
rect 23212 20728 23252 20768
rect 23116 20224 23156 20264
rect 25420 23836 25460 23876
rect 24556 23080 24596 23120
rect 26572 22324 26612 22364
rect 24172 22156 24212 22196
rect 23980 21484 24020 21524
rect 24172 21484 24212 21524
rect 23500 20140 23540 20180
rect 22732 19888 22772 19928
rect 23308 19888 23348 19928
rect 23500 19216 23540 19256
rect 22732 18460 22772 18500
rect 22636 18292 22676 18332
rect 22252 17620 22292 17660
rect 22252 17032 22292 17072
rect 22732 17704 22772 17744
rect 22924 17704 22964 17744
rect 22828 17620 22868 17660
rect 22540 17032 22580 17072
rect 23020 16948 23060 16988
rect 19472 14344 19512 14384
rect 19554 14344 19594 14384
rect 19636 14344 19676 14384
rect 19718 14344 19758 14384
rect 19800 14344 19840 14384
rect 19472 12832 19512 12872
rect 19554 12832 19594 12872
rect 19636 12832 19676 12872
rect 19718 12832 19758 12872
rect 19800 12832 19840 12872
rect 20140 12244 20180 12284
rect 26476 18712 26516 18752
rect 26092 18628 26132 18668
rect 26188 18460 26228 18500
rect 26380 18460 26420 18500
rect 26476 18292 26516 18332
rect 26284 17704 26324 17744
rect 26764 17704 26804 17744
rect 23788 15520 23828 15560
rect 25036 15520 25076 15560
rect 23020 12496 23060 12536
rect 26956 13168 26996 13208
rect 26860 12748 26900 12788
rect 26572 12664 26612 12704
rect 26476 12580 26516 12620
rect 26956 12664 26996 12704
rect 26764 12244 26804 12284
rect 24940 11908 24980 11948
rect 26380 11908 26420 11948
rect 19472 11320 19512 11360
rect 19554 11320 19594 11360
rect 19636 11320 19676 11360
rect 19718 11320 19758 11360
rect 19800 11320 19840 11360
rect 19472 9808 19512 9848
rect 19554 9808 19594 9848
rect 19636 9808 19676 9848
rect 19718 9808 19758 9848
rect 19800 9808 19840 9848
rect 27340 31144 27380 31184
rect 27148 28288 27188 28328
rect 27532 31900 27572 31940
rect 27916 31312 27956 31352
rect 28780 31228 28820 31268
rect 27628 30640 27668 30680
rect 28780 30556 28820 30596
rect 28300 30220 28340 30260
rect 28204 28456 28244 28496
rect 29164 30220 29204 30260
rect 28780 28456 28820 28496
rect 27532 28372 27572 28412
rect 28108 28288 28148 28328
rect 28012 28204 28052 28244
rect 28300 27784 28340 27824
rect 28108 27448 28148 27488
rect 28492 28120 28532 28160
rect 28396 27700 28436 27740
rect 34592 34000 34632 34040
rect 34674 34000 34714 34040
rect 34756 34000 34796 34040
rect 34838 34000 34878 34040
rect 34920 34000 34960 34040
rect 49712 34000 49752 34040
rect 49794 34000 49834 34040
rect 49876 34000 49916 34040
rect 49958 34000 49998 34040
rect 50040 34000 50080 34040
rect 64832 34000 64872 34040
rect 64914 34000 64954 34040
rect 64996 34000 65036 34040
rect 65078 34000 65118 34040
rect 65160 34000 65200 34040
rect 79952 34000 79992 34040
rect 80034 34000 80074 34040
rect 80116 34000 80156 34040
rect 80198 34000 80238 34040
rect 80280 34000 80320 34040
rect 95072 34000 95112 34040
rect 95154 34000 95194 34040
rect 95236 34000 95276 34040
rect 95318 34000 95358 34040
rect 95400 34000 95440 34040
rect 29644 33664 29684 33704
rect 33352 33244 33392 33284
rect 33434 33244 33474 33284
rect 33516 33244 33556 33284
rect 33598 33244 33638 33284
rect 33680 33244 33720 33284
rect 48472 33244 48512 33284
rect 48554 33244 48594 33284
rect 48636 33244 48676 33284
rect 48718 33244 48758 33284
rect 48800 33244 48840 33284
rect 63592 33244 63632 33284
rect 63674 33244 63714 33284
rect 63756 33244 63796 33284
rect 63838 33244 63878 33284
rect 63920 33244 63960 33284
rect 78712 33244 78752 33284
rect 78794 33244 78834 33284
rect 78876 33244 78916 33284
rect 78958 33244 78998 33284
rect 79040 33244 79080 33284
rect 93832 33244 93872 33284
rect 93914 33244 93954 33284
rect 93996 33244 94036 33284
rect 94078 33244 94118 33284
rect 94160 33244 94200 33284
rect 34592 32488 34632 32528
rect 34674 32488 34714 32528
rect 34756 32488 34796 32528
rect 34838 32488 34878 32528
rect 34920 32488 34960 32528
rect 49712 32488 49752 32528
rect 49794 32488 49834 32528
rect 49876 32488 49916 32528
rect 49958 32488 49998 32528
rect 50040 32488 50080 32528
rect 64832 32488 64872 32528
rect 64914 32488 64954 32528
rect 64996 32488 65036 32528
rect 65078 32488 65118 32528
rect 65160 32488 65200 32528
rect 79952 32488 79992 32528
rect 80034 32488 80074 32528
rect 80116 32488 80156 32528
rect 80198 32488 80238 32528
rect 80280 32488 80320 32528
rect 95072 32488 95112 32528
rect 95154 32488 95194 32528
rect 95236 32488 95276 32528
rect 95318 32488 95358 32528
rect 95400 32488 95440 32528
rect 33352 31732 33392 31772
rect 33434 31732 33474 31772
rect 33516 31732 33556 31772
rect 33598 31732 33638 31772
rect 33680 31732 33720 31772
rect 48472 31732 48512 31772
rect 48554 31732 48594 31772
rect 48636 31732 48676 31772
rect 48718 31732 48758 31772
rect 48800 31732 48840 31772
rect 63592 31732 63632 31772
rect 63674 31732 63714 31772
rect 63756 31732 63796 31772
rect 63838 31732 63878 31772
rect 63920 31732 63960 31772
rect 78712 31732 78752 31772
rect 78794 31732 78834 31772
rect 78876 31732 78916 31772
rect 78958 31732 78998 31772
rect 79040 31732 79080 31772
rect 93832 31732 93872 31772
rect 93914 31732 93954 31772
rect 93996 31732 94036 31772
rect 94078 31732 94118 31772
rect 94160 31732 94200 31772
rect 34592 30976 34632 31016
rect 34674 30976 34714 31016
rect 34756 30976 34796 31016
rect 34838 30976 34878 31016
rect 34920 30976 34960 31016
rect 49712 30976 49752 31016
rect 49794 30976 49834 31016
rect 49876 30976 49916 31016
rect 49958 30976 49998 31016
rect 50040 30976 50080 31016
rect 64832 30976 64872 31016
rect 64914 30976 64954 31016
rect 64996 30976 65036 31016
rect 65078 30976 65118 31016
rect 65160 30976 65200 31016
rect 79952 30976 79992 31016
rect 80034 30976 80074 31016
rect 80116 30976 80156 31016
rect 80198 30976 80238 31016
rect 80280 30976 80320 31016
rect 95072 30976 95112 31016
rect 95154 30976 95194 31016
rect 95236 30976 95276 31016
rect 95318 30976 95358 31016
rect 95400 30976 95440 31016
rect 32812 30640 32852 30680
rect 31276 30220 31316 30260
rect 32716 30220 32756 30260
rect 29452 28120 29492 28160
rect 29452 27700 29492 27740
rect 29164 27532 29204 27572
rect 29260 27448 29300 27488
rect 29452 27532 29492 27572
rect 29356 27364 29396 27404
rect 29644 27640 29684 27656
rect 29644 27616 29684 27640
rect 31180 28288 31220 28328
rect 30028 27532 30068 27572
rect 30124 27364 30164 27404
rect 28204 26020 28244 26060
rect 28204 25516 28244 25556
rect 28396 25264 28436 25304
rect 28012 25096 28052 25136
rect 28492 25096 28532 25136
rect 27532 24508 27572 24548
rect 29260 25264 29300 25304
rect 30028 25264 30068 25304
rect 28492 23668 28532 23708
rect 27244 22492 27284 22532
rect 28588 22828 28628 22868
rect 28972 23668 29012 23708
rect 28876 22576 28916 22616
rect 28684 22408 28724 22448
rect 28876 22408 28916 22448
rect 28780 22324 28820 22364
rect 28396 21568 28436 21608
rect 29164 22408 29204 22448
rect 29836 24508 29876 24548
rect 33964 30640 34004 30680
rect 33100 30556 33140 30596
rect 34348 30556 34388 30596
rect 33352 30220 33392 30260
rect 33434 30220 33474 30260
rect 33516 30220 33556 30260
rect 33598 30220 33638 30260
rect 33680 30220 33720 30260
rect 33352 28708 33392 28748
rect 33434 28708 33474 28748
rect 33516 28708 33556 28748
rect 33598 28708 33638 28748
rect 33680 28708 33720 28748
rect 33352 27196 33392 27236
rect 33434 27196 33474 27236
rect 33516 27196 33556 27236
rect 33598 27196 33638 27236
rect 33680 27196 33720 27236
rect 35116 30388 35156 30428
rect 35596 30388 35636 30428
rect 34592 29464 34632 29504
rect 34674 29464 34714 29504
rect 34756 29464 34796 29504
rect 34838 29464 34878 29504
rect 34920 29464 34960 29504
rect 48472 30220 48512 30260
rect 48554 30220 48594 30260
rect 48636 30220 48676 30260
rect 48718 30220 48758 30260
rect 48800 30220 48840 30260
rect 63592 30220 63632 30260
rect 63674 30220 63714 30260
rect 63756 30220 63796 30260
rect 63838 30220 63878 30260
rect 63920 30220 63960 30260
rect 78712 30220 78752 30260
rect 78794 30220 78834 30260
rect 78876 30220 78916 30260
rect 78958 30220 78998 30260
rect 79040 30220 79080 30260
rect 93832 30220 93872 30260
rect 93914 30220 93954 30260
rect 93996 30220 94036 30260
rect 94078 30220 94118 30260
rect 94160 30220 94200 30260
rect 34592 27952 34632 27992
rect 34674 27952 34714 27992
rect 34756 27952 34796 27992
rect 34838 27952 34878 27992
rect 34920 27952 34960 27992
rect 34924 27280 34964 27320
rect 35788 28960 35828 29000
rect 35884 27028 35924 27068
rect 34592 26440 34632 26480
rect 34674 26440 34714 26480
rect 34756 26440 34796 26480
rect 34838 26440 34878 26480
rect 34920 26440 34960 26480
rect 35404 26776 35444 26816
rect 35308 26020 35348 26060
rect 33352 25684 33392 25724
rect 33434 25684 33474 25724
rect 33516 25684 33556 25724
rect 33598 25684 33638 25724
rect 33680 25684 33720 25724
rect 35212 25180 35252 25220
rect 34592 24928 34632 24968
rect 34674 24928 34714 24968
rect 34756 24928 34796 24968
rect 34838 24928 34878 24968
rect 34920 24928 34960 24968
rect 35212 24508 35252 24548
rect 33352 24172 33392 24212
rect 33434 24172 33474 24212
rect 33516 24172 33556 24212
rect 33598 24172 33638 24212
rect 33680 24172 33720 24212
rect 32812 23836 32852 23876
rect 30124 23752 30164 23792
rect 29644 23668 29684 23708
rect 32812 23584 32852 23624
rect 32620 22492 32660 22532
rect 29164 20896 29204 20936
rect 28876 20812 28916 20852
rect 32524 22240 32564 22280
rect 32428 22072 32468 22112
rect 33100 21820 33140 21860
rect 29356 21568 29396 21608
rect 30316 20896 30356 20936
rect 29260 20728 29300 20768
rect 29644 20728 29684 20768
rect 31372 20812 31412 20852
rect 30508 20728 30548 20768
rect 28108 20140 28148 20180
rect 29452 20140 29492 20180
rect 27340 18628 27380 18668
rect 27436 18544 27476 18584
rect 28012 17704 28052 17744
rect 28396 18544 28436 18584
rect 28204 17620 28244 17660
rect 29164 17620 29204 17660
rect 27148 16948 27188 16988
rect 27916 15520 27956 15560
rect 30892 20560 30932 20600
rect 32620 18880 32660 18920
rect 31372 17788 31412 17828
rect 34444 23752 34484 23792
rect 33772 23584 33812 23624
rect 33352 22660 33392 22700
rect 33434 22660 33474 22700
rect 33516 22660 33556 22700
rect 33598 22660 33638 22700
rect 33680 22660 33720 22700
rect 34592 23416 34632 23456
rect 34674 23416 34714 23456
rect 34756 23416 34796 23456
rect 34838 23416 34878 23456
rect 34920 23416 34960 23456
rect 34156 22576 34196 22616
rect 34924 22576 34964 22616
rect 34060 22240 34100 22280
rect 34348 22324 34388 22364
rect 34732 22324 34772 22364
rect 34252 22156 34292 22196
rect 34156 22072 34196 22112
rect 33196 21568 33236 21608
rect 33352 21148 33392 21188
rect 33434 21148 33474 21188
rect 33516 21148 33556 21188
rect 33598 21148 33638 21188
rect 33680 21148 33720 21188
rect 34060 20644 34100 20684
rect 33772 20056 33812 20096
rect 33352 19636 33392 19676
rect 33434 19636 33474 19676
rect 33516 19636 33556 19676
rect 33598 19636 33638 19676
rect 33680 19636 33720 19676
rect 33352 18124 33392 18164
rect 33434 18124 33474 18164
rect 33516 18124 33556 18164
rect 33598 18124 33638 18164
rect 33680 18124 33720 18164
rect 33868 19216 33908 19256
rect 33868 18880 33908 18920
rect 32620 17704 32660 17744
rect 33100 17704 33140 17744
rect 31276 17032 31316 17072
rect 31756 17032 31796 17072
rect 31180 16948 31220 16988
rect 30604 16360 30644 16400
rect 28300 15436 28340 15476
rect 27820 12748 27860 12788
rect 27244 12580 27284 12620
rect 27436 12412 27476 12452
rect 28012 12412 28052 12452
rect 33676 17704 33716 17744
rect 33772 17620 33812 17660
rect 34060 16948 34100 16988
rect 33352 16612 33392 16652
rect 33434 16612 33474 16652
rect 33516 16612 33556 16652
rect 33598 16612 33638 16652
rect 33680 16612 33720 16652
rect 33196 16360 33236 16400
rect 33772 16360 33812 16400
rect 33100 15520 33140 15560
rect 34060 16276 34100 16316
rect 34348 21904 34388 21944
rect 34252 17620 34292 17660
rect 33352 15100 33392 15140
rect 33434 15100 33474 15140
rect 33516 15100 33556 15140
rect 33598 15100 33638 15140
rect 33680 15100 33720 15140
rect 33352 13588 33392 13628
rect 33434 13588 33474 13628
rect 33516 13588 33556 13628
rect 33598 13588 33638 13628
rect 33680 13588 33720 13628
rect 33196 13168 33236 13208
rect 33004 13000 33044 13040
rect 34156 13168 34196 13208
rect 27244 12244 27284 12284
rect 33352 12076 33392 12116
rect 33434 12076 33474 12116
rect 33516 12076 33556 12116
rect 33598 12076 33638 12116
rect 33680 12076 33720 12116
rect 27820 11992 27860 12032
rect 33352 10564 33392 10604
rect 33434 10564 33474 10604
rect 33516 10564 33556 10604
rect 33598 10564 33638 10604
rect 33680 10564 33720 10604
rect 27052 9388 27092 9428
rect 33352 9052 33392 9092
rect 33434 9052 33474 9092
rect 33516 9052 33556 9092
rect 33598 9052 33638 9092
rect 33680 9052 33720 9092
rect 19472 8296 19512 8336
rect 19554 8296 19594 8336
rect 19636 8296 19676 8336
rect 19718 8296 19758 8336
rect 19800 8296 19840 8336
rect 33352 7540 33392 7580
rect 33434 7540 33474 7580
rect 33516 7540 33556 7580
rect 33598 7540 33638 7580
rect 33680 7540 33720 7580
rect 34252 7204 34292 7244
rect 19472 6784 19512 6824
rect 19554 6784 19594 6824
rect 19636 6784 19676 6824
rect 19718 6784 19758 6824
rect 19800 6784 19840 6824
rect 3112 6028 3152 6068
rect 3194 6028 3234 6068
rect 3276 6028 3316 6068
rect 3358 6028 3398 6068
rect 3440 6028 3480 6068
rect 18232 6028 18272 6068
rect 18314 6028 18354 6068
rect 18396 6028 18436 6068
rect 18478 6028 18518 6068
rect 18560 6028 18600 6068
rect 33352 6028 33392 6068
rect 33434 6028 33474 6068
rect 33516 6028 33556 6068
rect 33598 6028 33638 6068
rect 33680 6028 33720 6068
rect 18700 5692 18740 5732
rect 4352 5272 4392 5312
rect 4434 5272 4474 5312
rect 4516 5272 4556 5312
rect 4598 5272 4638 5312
rect 4680 5272 4720 5312
rect 19472 5272 19512 5312
rect 19554 5272 19594 5312
rect 19636 5272 19676 5312
rect 19718 5272 19758 5312
rect 19800 5272 19840 5312
rect 34348 4852 34388 4892
rect 3112 4516 3152 4556
rect 3194 4516 3234 4556
rect 3276 4516 3316 4556
rect 3358 4516 3398 4556
rect 3440 4516 3480 4556
rect 18232 4516 18272 4556
rect 18314 4516 18354 4556
rect 18396 4516 18436 4556
rect 18478 4516 18518 4556
rect 18560 4516 18600 4556
rect 33352 4516 33392 4556
rect 33434 4516 33474 4556
rect 33516 4516 33556 4556
rect 33598 4516 33638 4556
rect 33680 4516 33720 4556
rect 34636 22072 34676 22112
rect 35500 26020 35540 26060
rect 35596 25180 35636 25220
rect 36460 28960 36500 29000
rect 36172 26776 36212 26816
rect 35500 23836 35540 23876
rect 35404 23584 35444 23624
rect 35308 23080 35348 23120
rect 35596 22408 35636 22448
rect 35980 22408 36020 22448
rect 35308 22324 35348 22364
rect 35020 22156 35060 22196
rect 34828 22072 34868 22112
rect 35020 21988 35060 22028
rect 34592 21904 34632 21944
rect 34674 21904 34714 21944
rect 34756 21904 34796 21944
rect 34838 21904 34878 21944
rect 34920 21904 34960 21944
rect 34592 20392 34632 20432
rect 34674 20392 34714 20432
rect 34756 20392 34796 20432
rect 34838 20392 34878 20432
rect 34920 20392 34960 20432
rect 35404 22240 35444 22280
rect 35788 22324 35828 22364
rect 36460 22240 36500 22280
rect 35692 22156 35732 22196
rect 35212 21820 35252 21860
rect 34828 20056 34868 20096
rect 35020 20056 35060 20096
rect 34592 18880 34632 18920
rect 34674 18880 34714 18920
rect 34756 18880 34796 18920
rect 34838 18880 34878 18920
rect 34920 18880 34960 18920
rect 34592 17368 34632 17408
rect 34674 17368 34714 17408
rect 34756 17368 34796 17408
rect 34838 17368 34878 17408
rect 34920 17368 34960 17408
rect 34592 15856 34632 15896
rect 34674 15856 34714 15896
rect 34756 15856 34796 15896
rect 34838 15856 34878 15896
rect 34920 15856 34960 15896
rect 34592 14344 34632 14384
rect 34674 14344 34714 14384
rect 34756 14344 34796 14384
rect 34838 14344 34878 14384
rect 34920 14344 34960 14384
rect 34592 12832 34632 12872
rect 34674 12832 34714 12872
rect 34756 12832 34796 12872
rect 34838 12832 34878 12872
rect 34920 12832 34960 12872
rect 34592 11320 34632 11360
rect 34674 11320 34714 11360
rect 34756 11320 34796 11360
rect 34838 11320 34878 11360
rect 34920 11320 34960 11360
rect 49712 29464 49752 29504
rect 49794 29464 49834 29504
rect 49876 29464 49916 29504
rect 49958 29464 49998 29504
rect 50040 29464 50080 29504
rect 64832 29464 64872 29504
rect 64914 29464 64954 29504
rect 64996 29464 65036 29504
rect 65078 29464 65118 29504
rect 65160 29464 65200 29504
rect 79952 29464 79992 29504
rect 80034 29464 80074 29504
rect 80116 29464 80156 29504
rect 80198 29464 80238 29504
rect 80280 29464 80320 29504
rect 95072 29464 95112 29504
rect 95154 29464 95194 29504
rect 95236 29464 95276 29504
rect 95318 29464 95358 29504
rect 95400 29464 95440 29504
rect 48472 28708 48512 28748
rect 48554 28708 48594 28748
rect 48636 28708 48676 28748
rect 48718 28708 48758 28748
rect 48800 28708 48840 28748
rect 63592 28708 63632 28748
rect 63674 28708 63714 28748
rect 63756 28708 63796 28748
rect 63838 28708 63878 28748
rect 63920 28708 63960 28748
rect 78712 28708 78752 28748
rect 78794 28708 78834 28748
rect 78876 28708 78916 28748
rect 78958 28708 78998 28748
rect 79040 28708 79080 28748
rect 93832 28708 93872 28748
rect 93914 28708 93954 28748
rect 93996 28708 94036 28748
rect 94078 28708 94118 28748
rect 94160 28708 94200 28748
rect 49712 27952 49752 27992
rect 49794 27952 49834 27992
rect 49876 27952 49916 27992
rect 49958 27952 49998 27992
rect 50040 27952 50080 27992
rect 64832 27952 64872 27992
rect 64914 27952 64954 27992
rect 64996 27952 65036 27992
rect 65078 27952 65118 27992
rect 65160 27952 65200 27992
rect 79952 27952 79992 27992
rect 80034 27952 80074 27992
rect 80116 27952 80156 27992
rect 80198 27952 80238 27992
rect 80280 27952 80320 27992
rect 95072 27952 95112 27992
rect 95154 27952 95194 27992
rect 95236 27952 95276 27992
rect 95318 27952 95358 27992
rect 95400 27952 95440 27992
rect 48472 27196 48512 27236
rect 48554 27196 48594 27236
rect 48636 27196 48676 27236
rect 48718 27196 48758 27236
rect 48800 27196 48840 27236
rect 63592 27196 63632 27236
rect 63674 27196 63714 27236
rect 63756 27196 63796 27236
rect 63838 27196 63878 27236
rect 63920 27196 63960 27236
rect 78712 27196 78752 27236
rect 78794 27196 78834 27236
rect 78876 27196 78916 27236
rect 78958 27196 78998 27236
rect 79040 27196 79080 27236
rect 93832 27196 93872 27236
rect 93914 27196 93954 27236
rect 93996 27196 94036 27236
rect 94078 27196 94118 27236
rect 94160 27196 94200 27236
rect 37324 27028 37364 27068
rect 49712 26440 49752 26480
rect 49794 26440 49834 26480
rect 49876 26440 49916 26480
rect 49958 26440 49998 26480
rect 50040 26440 50080 26480
rect 64832 26440 64872 26480
rect 64914 26440 64954 26480
rect 64996 26440 65036 26480
rect 65078 26440 65118 26480
rect 65160 26440 65200 26480
rect 79952 26440 79992 26480
rect 80034 26440 80074 26480
rect 80116 26440 80156 26480
rect 80198 26440 80238 26480
rect 80280 26440 80320 26480
rect 95072 26440 95112 26480
rect 95154 26440 95194 26480
rect 95236 26440 95276 26480
rect 95318 26440 95358 26480
rect 95400 26440 95440 26480
rect 39628 26104 39668 26144
rect 48472 25684 48512 25724
rect 48554 25684 48594 25724
rect 48636 25684 48676 25724
rect 48718 25684 48758 25724
rect 48800 25684 48840 25724
rect 63592 25684 63632 25724
rect 63674 25684 63714 25724
rect 63756 25684 63796 25724
rect 63838 25684 63878 25724
rect 63920 25684 63960 25724
rect 78712 25684 78752 25724
rect 78794 25684 78834 25724
rect 78876 25684 78916 25724
rect 78958 25684 78998 25724
rect 79040 25684 79080 25724
rect 93832 25684 93872 25724
rect 93914 25684 93954 25724
rect 93996 25684 94036 25724
rect 94078 25684 94118 25724
rect 94160 25684 94200 25724
rect 49712 24928 49752 24968
rect 49794 24928 49834 24968
rect 49876 24928 49916 24968
rect 49958 24928 49998 24968
rect 50040 24928 50080 24968
rect 64832 24928 64872 24968
rect 64914 24928 64954 24968
rect 64996 24928 65036 24968
rect 65078 24928 65118 24968
rect 65160 24928 65200 24968
rect 79952 24928 79992 24968
rect 80034 24928 80074 24968
rect 80116 24928 80156 24968
rect 80198 24928 80238 24968
rect 80280 24928 80320 24968
rect 95072 24928 95112 24968
rect 95154 24928 95194 24968
rect 95236 24928 95276 24968
rect 95318 24928 95358 24968
rect 95400 24928 95440 24968
rect 48472 24172 48512 24212
rect 48554 24172 48594 24212
rect 48636 24172 48676 24212
rect 48718 24172 48758 24212
rect 48800 24172 48840 24212
rect 63592 24172 63632 24212
rect 63674 24172 63714 24212
rect 63756 24172 63796 24212
rect 63838 24172 63878 24212
rect 63920 24172 63960 24212
rect 78712 24172 78752 24212
rect 78794 24172 78834 24212
rect 78876 24172 78916 24212
rect 78958 24172 78998 24212
rect 79040 24172 79080 24212
rect 93832 24172 93872 24212
rect 93914 24172 93954 24212
rect 93996 24172 94036 24212
rect 94078 24172 94118 24212
rect 94160 24172 94200 24212
rect 39916 23836 39956 23876
rect 49712 23416 49752 23456
rect 49794 23416 49834 23456
rect 49876 23416 49916 23456
rect 49958 23416 49998 23456
rect 50040 23416 50080 23456
rect 64832 23416 64872 23456
rect 64914 23416 64954 23456
rect 64996 23416 65036 23456
rect 65078 23416 65118 23456
rect 65160 23416 65200 23456
rect 79952 23416 79992 23456
rect 80034 23416 80074 23456
rect 80116 23416 80156 23456
rect 80198 23416 80238 23456
rect 80280 23416 80320 23456
rect 95072 23416 95112 23456
rect 95154 23416 95194 23456
rect 95236 23416 95276 23456
rect 95318 23416 95358 23456
rect 95400 23416 95440 23456
rect 40396 23080 40436 23120
rect 39532 22660 39572 22700
rect 39916 22660 39956 22700
rect 37228 19804 37268 19844
rect 37036 19300 37076 19340
rect 37516 19384 37556 19424
rect 38764 19384 38804 19424
rect 38860 19216 38900 19256
rect 38764 19048 38804 19088
rect 36844 18628 36884 18668
rect 37228 18628 37268 18668
rect 37900 17116 37940 17156
rect 37324 16192 37364 16232
rect 38572 16192 38612 16232
rect 39244 19804 39284 19844
rect 48472 22660 48512 22700
rect 48554 22660 48594 22700
rect 48636 22660 48676 22700
rect 48718 22660 48758 22700
rect 48800 22660 48840 22700
rect 63592 22660 63632 22700
rect 63674 22660 63714 22700
rect 63756 22660 63796 22700
rect 63838 22660 63878 22700
rect 63920 22660 63960 22700
rect 78712 22660 78752 22700
rect 78794 22660 78834 22700
rect 78876 22660 78916 22700
rect 78958 22660 78998 22700
rect 79040 22660 79080 22700
rect 93832 22660 93872 22700
rect 93914 22660 93954 22700
rect 93996 22660 94036 22700
rect 94078 22660 94118 22700
rect 94160 22660 94200 22700
rect 41548 22324 41588 22364
rect 49712 21904 49752 21944
rect 49794 21904 49834 21944
rect 49876 21904 49916 21944
rect 49958 21904 49998 21944
rect 50040 21904 50080 21944
rect 64832 21904 64872 21944
rect 64914 21904 64954 21944
rect 64996 21904 65036 21944
rect 65078 21904 65118 21944
rect 65160 21904 65200 21944
rect 79952 21904 79992 21944
rect 80034 21904 80074 21944
rect 80116 21904 80156 21944
rect 80198 21904 80238 21944
rect 80280 21904 80320 21944
rect 95072 21904 95112 21944
rect 95154 21904 95194 21944
rect 95236 21904 95276 21944
rect 95318 21904 95358 21944
rect 95400 21904 95440 21944
rect 48472 21148 48512 21188
rect 48554 21148 48594 21188
rect 48636 21148 48676 21188
rect 48718 21148 48758 21188
rect 48800 21148 48840 21188
rect 63592 21148 63632 21188
rect 63674 21148 63714 21188
rect 63756 21148 63796 21188
rect 63838 21148 63878 21188
rect 63920 21148 63960 21188
rect 78712 21148 78752 21188
rect 78794 21148 78834 21188
rect 78876 21148 78916 21188
rect 78958 21148 78998 21188
rect 79040 21148 79080 21188
rect 93832 21148 93872 21188
rect 93914 21148 93954 21188
rect 93996 21148 94036 21188
rect 94078 21148 94118 21188
rect 94160 21148 94200 21188
rect 49712 20392 49752 20432
rect 49794 20392 49834 20432
rect 49876 20392 49916 20432
rect 49958 20392 49998 20432
rect 50040 20392 50080 20432
rect 64832 20392 64872 20432
rect 64914 20392 64954 20432
rect 64996 20392 65036 20432
rect 65078 20392 65118 20432
rect 65160 20392 65200 20432
rect 79952 20392 79992 20432
rect 80034 20392 80074 20432
rect 80116 20392 80156 20432
rect 80198 20392 80238 20432
rect 80280 20392 80320 20432
rect 95072 20392 95112 20432
rect 95154 20392 95194 20432
rect 95236 20392 95276 20432
rect 95318 20392 95358 20432
rect 95400 20392 95440 20432
rect 39916 20056 39956 20096
rect 41164 20056 41204 20096
rect 48472 19636 48512 19676
rect 48554 19636 48594 19676
rect 48636 19636 48676 19676
rect 48718 19636 48758 19676
rect 48800 19636 48840 19676
rect 63592 19636 63632 19676
rect 63674 19636 63714 19676
rect 63756 19636 63796 19676
rect 63838 19636 63878 19676
rect 63920 19636 63960 19676
rect 78712 19636 78752 19676
rect 78794 19636 78834 19676
rect 78876 19636 78916 19676
rect 78958 19636 78998 19676
rect 79040 19636 79080 19676
rect 93832 19636 93872 19676
rect 93914 19636 93954 19676
rect 93996 19636 94036 19676
rect 94078 19636 94118 19676
rect 94160 19636 94200 19676
rect 40012 19216 40052 19256
rect 39148 19048 39188 19088
rect 39532 19048 39572 19088
rect 49712 18880 49752 18920
rect 49794 18880 49834 18920
rect 49876 18880 49916 18920
rect 49958 18880 49998 18920
rect 50040 18880 50080 18920
rect 64832 18880 64872 18920
rect 64914 18880 64954 18920
rect 64996 18880 65036 18920
rect 65078 18880 65118 18920
rect 65160 18880 65200 18920
rect 79952 18880 79992 18920
rect 80034 18880 80074 18920
rect 80116 18880 80156 18920
rect 80198 18880 80238 18920
rect 80280 18880 80320 18920
rect 95072 18880 95112 18920
rect 95154 18880 95194 18920
rect 95236 18880 95276 18920
rect 95318 18880 95358 18920
rect 95400 18880 95440 18920
rect 39052 18460 39092 18500
rect 48472 18124 48512 18164
rect 48554 18124 48594 18164
rect 48636 18124 48676 18164
rect 48718 18124 48758 18164
rect 48800 18124 48840 18164
rect 63592 18124 63632 18164
rect 63674 18124 63714 18164
rect 63756 18124 63796 18164
rect 63838 18124 63878 18164
rect 63920 18124 63960 18164
rect 78712 18124 78752 18164
rect 78794 18124 78834 18164
rect 78876 18124 78916 18164
rect 78958 18124 78998 18164
rect 79040 18124 79080 18164
rect 93832 18124 93872 18164
rect 93914 18124 93954 18164
rect 93996 18124 94036 18164
rect 94078 18124 94118 18164
rect 94160 18124 94200 18164
rect 49712 17368 49752 17408
rect 49794 17368 49834 17408
rect 49876 17368 49916 17408
rect 49958 17368 49998 17408
rect 50040 17368 50080 17408
rect 64832 17368 64872 17408
rect 64914 17368 64954 17408
rect 64996 17368 65036 17408
rect 65078 17368 65118 17408
rect 65160 17368 65200 17408
rect 79952 17368 79992 17408
rect 80034 17368 80074 17408
rect 80116 17368 80156 17408
rect 80198 17368 80238 17408
rect 80280 17368 80320 17408
rect 95072 17368 95112 17408
rect 95154 17368 95194 17408
rect 95236 17368 95276 17408
rect 95318 17368 95358 17408
rect 95400 17368 95440 17408
rect 48472 16612 48512 16652
rect 48554 16612 48594 16652
rect 48636 16612 48676 16652
rect 48718 16612 48758 16652
rect 48800 16612 48840 16652
rect 63592 16612 63632 16652
rect 63674 16612 63714 16652
rect 63756 16612 63796 16652
rect 63838 16612 63878 16652
rect 63920 16612 63960 16652
rect 78712 16612 78752 16652
rect 78794 16612 78834 16652
rect 78876 16612 78916 16652
rect 78958 16612 78998 16652
rect 79040 16612 79080 16652
rect 93832 16612 93872 16652
rect 93914 16612 93954 16652
rect 93996 16612 94036 16652
rect 94078 16612 94118 16652
rect 94160 16612 94200 16652
rect 39244 16276 39284 16316
rect 40012 16276 40052 16316
rect 49712 15856 49752 15896
rect 49794 15856 49834 15896
rect 49876 15856 49916 15896
rect 49958 15856 49998 15896
rect 50040 15856 50080 15896
rect 64832 15856 64872 15896
rect 64914 15856 64954 15896
rect 64996 15856 65036 15896
rect 65078 15856 65118 15896
rect 65160 15856 65200 15896
rect 79952 15856 79992 15896
rect 80034 15856 80074 15896
rect 80116 15856 80156 15896
rect 80198 15856 80238 15896
rect 80280 15856 80320 15896
rect 95072 15856 95112 15896
rect 95154 15856 95194 15896
rect 95236 15856 95276 15896
rect 95318 15856 95358 15896
rect 95400 15856 95440 15896
rect 48472 15100 48512 15140
rect 48554 15100 48594 15140
rect 48636 15100 48676 15140
rect 48718 15100 48758 15140
rect 48800 15100 48840 15140
rect 63592 15100 63632 15140
rect 63674 15100 63714 15140
rect 63756 15100 63796 15140
rect 63838 15100 63878 15140
rect 63920 15100 63960 15140
rect 78712 15100 78752 15140
rect 78794 15100 78834 15140
rect 78876 15100 78916 15140
rect 78958 15100 78998 15140
rect 79040 15100 79080 15140
rect 93832 15100 93872 15140
rect 93914 15100 93954 15140
rect 93996 15100 94036 15140
rect 94078 15100 94118 15140
rect 94160 15100 94200 15140
rect 49712 14344 49752 14384
rect 49794 14344 49834 14384
rect 49876 14344 49916 14384
rect 49958 14344 49998 14384
rect 50040 14344 50080 14384
rect 64832 14344 64872 14384
rect 64914 14344 64954 14384
rect 64996 14344 65036 14384
rect 65078 14344 65118 14384
rect 65160 14344 65200 14384
rect 79952 14344 79992 14384
rect 80034 14344 80074 14384
rect 80116 14344 80156 14384
rect 80198 14344 80238 14384
rect 80280 14344 80320 14384
rect 95072 14344 95112 14384
rect 95154 14344 95194 14384
rect 95236 14344 95276 14384
rect 95318 14344 95358 14384
rect 95400 14344 95440 14384
rect 48472 13588 48512 13628
rect 48554 13588 48594 13628
rect 48636 13588 48676 13628
rect 48718 13588 48758 13628
rect 48800 13588 48840 13628
rect 63592 13588 63632 13628
rect 63674 13588 63714 13628
rect 63756 13588 63796 13628
rect 63838 13588 63878 13628
rect 63920 13588 63960 13628
rect 78712 13588 78752 13628
rect 78794 13588 78834 13628
rect 78876 13588 78916 13628
rect 78958 13588 78998 13628
rect 79040 13588 79080 13628
rect 93832 13588 93872 13628
rect 93914 13588 93954 13628
rect 93996 13588 94036 13628
rect 94078 13588 94118 13628
rect 94160 13588 94200 13628
rect 49712 12832 49752 12872
rect 49794 12832 49834 12872
rect 49876 12832 49916 12872
rect 49958 12832 49998 12872
rect 50040 12832 50080 12872
rect 64832 12832 64872 12872
rect 64914 12832 64954 12872
rect 64996 12832 65036 12872
rect 65078 12832 65118 12872
rect 65160 12832 65200 12872
rect 79952 12832 79992 12872
rect 80034 12832 80074 12872
rect 80116 12832 80156 12872
rect 80198 12832 80238 12872
rect 80280 12832 80320 12872
rect 95072 12832 95112 12872
rect 95154 12832 95194 12872
rect 95236 12832 95276 12872
rect 95318 12832 95358 12872
rect 95400 12832 95440 12872
rect 48472 12076 48512 12116
rect 48554 12076 48594 12116
rect 48636 12076 48676 12116
rect 48718 12076 48758 12116
rect 48800 12076 48840 12116
rect 63592 12076 63632 12116
rect 63674 12076 63714 12116
rect 63756 12076 63796 12116
rect 63838 12076 63878 12116
rect 63920 12076 63960 12116
rect 78712 12076 78752 12116
rect 78794 12076 78834 12116
rect 78876 12076 78916 12116
rect 78958 12076 78998 12116
rect 79040 12076 79080 12116
rect 93832 12076 93872 12116
rect 93914 12076 93954 12116
rect 93996 12076 94036 12116
rect 94078 12076 94118 12116
rect 94160 12076 94200 12116
rect 49712 11320 49752 11360
rect 49794 11320 49834 11360
rect 49876 11320 49916 11360
rect 49958 11320 49998 11360
rect 50040 11320 50080 11360
rect 64832 11320 64872 11360
rect 64914 11320 64954 11360
rect 64996 11320 65036 11360
rect 65078 11320 65118 11360
rect 65160 11320 65200 11360
rect 79952 11320 79992 11360
rect 80034 11320 80074 11360
rect 80116 11320 80156 11360
rect 80198 11320 80238 11360
rect 80280 11320 80320 11360
rect 95072 11320 95112 11360
rect 95154 11320 95194 11360
rect 95236 11320 95276 11360
rect 95318 11320 95358 11360
rect 95400 11320 95440 11360
rect 48472 10564 48512 10604
rect 48554 10564 48594 10604
rect 48636 10564 48676 10604
rect 48718 10564 48758 10604
rect 48800 10564 48840 10604
rect 63592 10564 63632 10604
rect 63674 10564 63714 10604
rect 63756 10564 63796 10604
rect 63838 10564 63878 10604
rect 63920 10564 63960 10604
rect 78712 10564 78752 10604
rect 78794 10564 78834 10604
rect 78876 10564 78916 10604
rect 78958 10564 78998 10604
rect 79040 10564 79080 10604
rect 93832 10564 93872 10604
rect 93914 10564 93954 10604
rect 93996 10564 94036 10604
rect 94078 10564 94118 10604
rect 94160 10564 94200 10604
rect 36748 10228 36788 10268
rect 34592 9808 34632 9848
rect 34674 9808 34714 9848
rect 34756 9808 34796 9848
rect 34838 9808 34878 9848
rect 34920 9808 34960 9848
rect 49712 9808 49752 9848
rect 49794 9808 49834 9848
rect 49876 9808 49916 9848
rect 49958 9808 49998 9848
rect 50040 9808 50080 9848
rect 64832 9808 64872 9848
rect 64914 9808 64954 9848
rect 64996 9808 65036 9848
rect 65078 9808 65118 9848
rect 65160 9808 65200 9848
rect 79952 9808 79992 9848
rect 80034 9808 80074 9848
rect 80116 9808 80156 9848
rect 80198 9808 80238 9848
rect 80280 9808 80320 9848
rect 95072 9808 95112 9848
rect 95154 9808 95194 9848
rect 95236 9808 95276 9848
rect 95318 9808 95358 9848
rect 95400 9808 95440 9848
rect 48472 9052 48512 9092
rect 48554 9052 48594 9092
rect 48636 9052 48676 9092
rect 48718 9052 48758 9092
rect 48800 9052 48840 9092
rect 63592 9052 63632 9092
rect 63674 9052 63714 9092
rect 63756 9052 63796 9092
rect 63838 9052 63878 9092
rect 63920 9052 63960 9092
rect 78712 9052 78752 9092
rect 78794 9052 78834 9092
rect 78876 9052 78916 9092
rect 78958 9052 78998 9092
rect 79040 9052 79080 9092
rect 93832 9052 93872 9092
rect 93914 9052 93954 9092
rect 93996 9052 94036 9092
rect 94078 9052 94118 9092
rect 94160 9052 94200 9092
rect 34592 8296 34632 8336
rect 34674 8296 34714 8336
rect 34756 8296 34796 8336
rect 34838 8296 34878 8336
rect 34920 8296 34960 8336
rect 49712 8296 49752 8336
rect 49794 8296 49834 8336
rect 49876 8296 49916 8336
rect 49958 8296 49998 8336
rect 50040 8296 50080 8336
rect 64832 8296 64872 8336
rect 64914 8296 64954 8336
rect 64996 8296 65036 8336
rect 65078 8296 65118 8336
rect 65160 8296 65200 8336
rect 79952 8296 79992 8336
rect 80034 8296 80074 8336
rect 80116 8296 80156 8336
rect 80198 8296 80238 8336
rect 80280 8296 80320 8336
rect 95072 8296 95112 8336
rect 95154 8296 95194 8336
rect 95236 8296 95276 8336
rect 95318 8296 95358 8336
rect 95400 8296 95440 8336
rect 48472 7540 48512 7580
rect 48554 7540 48594 7580
rect 48636 7540 48676 7580
rect 48718 7540 48758 7580
rect 48800 7540 48840 7580
rect 63592 7540 63632 7580
rect 63674 7540 63714 7580
rect 63756 7540 63796 7580
rect 63838 7540 63878 7580
rect 63920 7540 63960 7580
rect 78712 7540 78752 7580
rect 78794 7540 78834 7580
rect 78876 7540 78916 7580
rect 78958 7540 78998 7580
rect 79040 7540 79080 7580
rect 93832 7540 93872 7580
rect 93914 7540 93954 7580
rect 93996 7540 94036 7580
rect 94078 7540 94118 7580
rect 94160 7540 94200 7580
rect 34592 6784 34632 6824
rect 34674 6784 34714 6824
rect 34756 6784 34796 6824
rect 34838 6784 34878 6824
rect 34920 6784 34960 6824
rect 49712 6784 49752 6824
rect 49794 6784 49834 6824
rect 49876 6784 49916 6824
rect 49958 6784 49998 6824
rect 50040 6784 50080 6824
rect 64832 6784 64872 6824
rect 64914 6784 64954 6824
rect 64996 6784 65036 6824
rect 65078 6784 65118 6824
rect 65160 6784 65200 6824
rect 79952 6784 79992 6824
rect 80034 6784 80074 6824
rect 80116 6784 80156 6824
rect 80198 6784 80238 6824
rect 80280 6784 80320 6824
rect 95072 6784 95112 6824
rect 95154 6784 95194 6824
rect 95236 6784 95276 6824
rect 95318 6784 95358 6824
rect 95400 6784 95440 6824
rect 48472 6028 48512 6068
rect 48554 6028 48594 6068
rect 48636 6028 48676 6068
rect 48718 6028 48758 6068
rect 48800 6028 48840 6068
rect 63592 6028 63632 6068
rect 63674 6028 63714 6068
rect 63756 6028 63796 6068
rect 63838 6028 63878 6068
rect 63920 6028 63960 6068
rect 78712 6028 78752 6068
rect 78794 6028 78834 6068
rect 78876 6028 78916 6068
rect 78958 6028 78998 6068
rect 79040 6028 79080 6068
rect 93832 6028 93872 6068
rect 93914 6028 93954 6068
rect 93996 6028 94036 6068
rect 94078 6028 94118 6068
rect 94160 6028 94200 6068
rect 34592 5272 34632 5312
rect 34674 5272 34714 5312
rect 34756 5272 34796 5312
rect 34838 5272 34878 5312
rect 34920 5272 34960 5312
rect 49712 5272 49752 5312
rect 49794 5272 49834 5312
rect 49876 5272 49916 5312
rect 49958 5272 49998 5312
rect 50040 5272 50080 5312
rect 64832 5272 64872 5312
rect 64914 5272 64954 5312
rect 64996 5272 65036 5312
rect 65078 5272 65118 5312
rect 65160 5272 65200 5312
rect 79952 5272 79992 5312
rect 80034 5272 80074 5312
rect 80116 5272 80156 5312
rect 80198 5272 80238 5312
rect 80280 5272 80320 5312
rect 95072 5272 95112 5312
rect 95154 5272 95194 5312
rect 95236 5272 95276 5312
rect 95318 5272 95358 5312
rect 95400 5272 95440 5312
rect 48472 4516 48512 4556
rect 48554 4516 48594 4556
rect 48636 4516 48676 4556
rect 48718 4516 48758 4556
rect 48800 4516 48840 4556
rect 63592 4516 63632 4556
rect 63674 4516 63714 4556
rect 63756 4516 63796 4556
rect 63838 4516 63878 4556
rect 63920 4516 63960 4556
rect 78712 4516 78752 4556
rect 78794 4516 78834 4556
rect 78876 4516 78916 4556
rect 78958 4516 78998 4556
rect 79040 4516 79080 4556
rect 93832 4516 93872 4556
rect 93914 4516 93954 4556
rect 93996 4516 94036 4556
rect 94078 4516 94118 4556
rect 94160 4516 94200 4556
rect 34444 4180 34484 4220
rect 4352 3760 4392 3800
rect 4434 3760 4474 3800
rect 4516 3760 4556 3800
rect 4598 3760 4638 3800
rect 4680 3760 4720 3800
rect 19472 3760 19512 3800
rect 19554 3760 19594 3800
rect 19636 3760 19676 3800
rect 19718 3760 19758 3800
rect 19800 3760 19840 3800
rect 34592 3760 34632 3800
rect 34674 3760 34714 3800
rect 34756 3760 34796 3800
rect 34838 3760 34878 3800
rect 34920 3760 34960 3800
rect 49712 3760 49752 3800
rect 49794 3760 49834 3800
rect 49876 3760 49916 3800
rect 49958 3760 49998 3800
rect 50040 3760 50080 3800
rect 64832 3760 64872 3800
rect 64914 3760 64954 3800
rect 64996 3760 65036 3800
rect 65078 3760 65118 3800
rect 65160 3760 65200 3800
rect 79952 3760 79992 3800
rect 80034 3760 80074 3800
rect 80116 3760 80156 3800
rect 80198 3760 80238 3800
rect 80280 3760 80320 3800
rect 95072 3760 95112 3800
rect 95154 3760 95194 3800
rect 95236 3760 95276 3800
rect 95318 3760 95358 3800
rect 95400 3760 95440 3800
rect 3112 3004 3152 3044
rect 3194 3004 3234 3044
rect 3276 3004 3316 3044
rect 3358 3004 3398 3044
rect 3440 3004 3480 3044
rect 18232 3004 18272 3044
rect 18314 3004 18354 3044
rect 18396 3004 18436 3044
rect 18478 3004 18518 3044
rect 18560 3004 18600 3044
rect 33352 3004 33392 3044
rect 33434 3004 33474 3044
rect 33516 3004 33556 3044
rect 33598 3004 33638 3044
rect 33680 3004 33720 3044
rect 48472 3004 48512 3044
rect 48554 3004 48594 3044
rect 48636 3004 48676 3044
rect 48718 3004 48758 3044
rect 48800 3004 48840 3044
rect 63592 3004 63632 3044
rect 63674 3004 63714 3044
rect 63756 3004 63796 3044
rect 63838 3004 63878 3044
rect 63920 3004 63960 3044
rect 78712 3004 78752 3044
rect 78794 3004 78834 3044
rect 78876 3004 78916 3044
rect 78958 3004 78998 3044
rect 79040 3004 79080 3044
rect 93832 3004 93872 3044
rect 93914 3004 93954 3044
rect 93996 3004 94036 3044
rect 94078 3004 94118 3044
rect 94160 3004 94200 3044
rect 652 2248 692 2288
rect 4352 2248 4392 2288
rect 4434 2248 4474 2288
rect 4516 2248 4556 2288
rect 4598 2248 4638 2288
rect 4680 2248 4720 2288
rect 19472 2248 19512 2288
rect 19554 2248 19594 2288
rect 19636 2248 19676 2288
rect 19718 2248 19758 2288
rect 19800 2248 19840 2288
rect 34592 2248 34632 2288
rect 34674 2248 34714 2288
rect 34756 2248 34796 2288
rect 34838 2248 34878 2288
rect 34920 2248 34960 2288
rect 49712 2248 49752 2288
rect 49794 2248 49834 2288
rect 49876 2248 49916 2288
rect 49958 2248 49998 2288
rect 50040 2248 50080 2288
rect 64832 2248 64872 2288
rect 64914 2248 64954 2288
rect 64996 2248 65036 2288
rect 65078 2248 65118 2288
rect 65160 2248 65200 2288
rect 79952 2248 79992 2288
rect 80034 2248 80074 2288
rect 80116 2248 80156 2288
rect 80198 2248 80238 2288
rect 80280 2248 80320 2288
rect 95072 2248 95112 2288
rect 95154 2248 95194 2288
rect 95236 2248 95276 2288
rect 95318 2248 95358 2288
rect 95400 2248 95440 2288
rect 3112 1492 3152 1532
rect 3194 1492 3234 1532
rect 3276 1492 3316 1532
rect 3358 1492 3398 1532
rect 3440 1492 3480 1532
rect 18232 1492 18272 1532
rect 18314 1492 18354 1532
rect 18396 1492 18436 1532
rect 18478 1492 18518 1532
rect 18560 1492 18600 1532
rect 33352 1492 33392 1532
rect 33434 1492 33474 1532
rect 33516 1492 33556 1532
rect 33598 1492 33638 1532
rect 33680 1492 33720 1532
rect 48472 1492 48512 1532
rect 48554 1492 48594 1532
rect 48636 1492 48676 1532
rect 48718 1492 48758 1532
rect 48800 1492 48840 1532
rect 63592 1492 63632 1532
rect 63674 1492 63714 1532
rect 63756 1492 63796 1532
rect 63838 1492 63878 1532
rect 63920 1492 63960 1532
rect 78712 1492 78752 1532
rect 78794 1492 78834 1532
rect 78876 1492 78916 1532
rect 78958 1492 78998 1532
rect 79040 1492 79080 1532
rect 93832 1492 93872 1532
rect 93914 1492 93954 1532
rect 93996 1492 94036 1532
rect 94078 1492 94118 1532
rect 94160 1492 94200 1532
rect 4352 736 4392 776
rect 4434 736 4474 776
rect 4516 736 4556 776
rect 4598 736 4638 776
rect 4680 736 4720 776
rect 19472 736 19512 776
rect 19554 736 19594 776
rect 19636 736 19676 776
rect 19718 736 19758 776
rect 19800 736 19840 776
rect 34592 736 34632 776
rect 34674 736 34714 776
rect 34756 736 34796 776
rect 34838 736 34878 776
rect 34920 736 34960 776
rect 49712 736 49752 776
rect 49794 736 49834 776
rect 49876 736 49916 776
rect 49958 736 49998 776
rect 50040 736 50080 776
rect 64832 736 64872 776
rect 64914 736 64954 776
rect 64996 736 65036 776
rect 65078 736 65118 776
rect 65160 736 65200 776
rect 79952 736 79992 776
rect 80034 736 80074 776
rect 80116 736 80156 776
rect 80198 736 80238 776
rect 80280 736 80320 776
rect 95072 736 95112 776
rect 95154 736 95194 776
rect 95236 736 95276 776
rect 95318 736 95358 776
rect 95400 736 95440 776
<< metal3 >>
rect 4343 38536 4352 38576
rect 4392 38536 4434 38576
rect 4474 38536 4516 38576
rect 4556 38536 4598 38576
rect 4638 38536 4680 38576
rect 4720 38536 4729 38576
rect 19463 38536 19472 38576
rect 19512 38536 19554 38576
rect 19594 38536 19636 38576
rect 19676 38536 19718 38576
rect 19758 38536 19800 38576
rect 19840 38536 19849 38576
rect 34583 38536 34592 38576
rect 34632 38536 34674 38576
rect 34714 38536 34756 38576
rect 34796 38536 34838 38576
rect 34878 38536 34920 38576
rect 34960 38536 34969 38576
rect 49703 38536 49712 38576
rect 49752 38536 49794 38576
rect 49834 38536 49876 38576
rect 49916 38536 49958 38576
rect 49998 38536 50040 38576
rect 50080 38536 50089 38576
rect 64823 38536 64832 38576
rect 64872 38536 64914 38576
rect 64954 38536 64996 38576
rect 65036 38536 65078 38576
rect 65118 38536 65160 38576
rect 65200 38536 65209 38576
rect 79943 38536 79952 38576
rect 79992 38536 80034 38576
rect 80074 38536 80116 38576
rect 80156 38536 80198 38576
rect 80238 38536 80280 38576
rect 80320 38536 80329 38576
rect 95063 38536 95072 38576
rect 95112 38536 95154 38576
rect 95194 38536 95236 38576
rect 95276 38536 95318 38576
rect 95358 38536 95400 38576
rect 95440 38536 95449 38576
rect 3103 37780 3112 37820
rect 3152 37780 3194 37820
rect 3234 37780 3276 37820
rect 3316 37780 3358 37820
rect 3398 37780 3440 37820
rect 3480 37780 3489 37820
rect 18223 37780 18232 37820
rect 18272 37780 18314 37820
rect 18354 37780 18396 37820
rect 18436 37780 18478 37820
rect 18518 37780 18560 37820
rect 18600 37780 18609 37820
rect 33343 37780 33352 37820
rect 33392 37780 33434 37820
rect 33474 37780 33516 37820
rect 33556 37780 33598 37820
rect 33638 37780 33680 37820
rect 33720 37780 33729 37820
rect 48463 37780 48472 37820
rect 48512 37780 48554 37820
rect 48594 37780 48636 37820
rect 48676 37780 48718 37820
rect 48758 37780 48800 37820
rect 48840 37780 48849 37820
rect 63583 37780 63592 37820
rect 63632 37780 63674 37820
rect 63714 37780 63756 37820
rect 63796 37780 63838 37820
rect 63878 37780 63920 37820
rect 63960 37780 63969 37820
rect 78703 37780 78712 37820
rect 78752 37780 78794 37820
rect 78834 37780 78876 37820
rect 78916 37780 78958 37820
rect 78998 37780 79040 37820
rect 79080 37780 79089 37820
rect 93823 37780 93832 37820
rect 93872 37780 93914 37820
rect 93954 37780 93996 37820
rect 94036 37780 94078 37820
rect 94118 37780 94160 37820
rect 94200 37780 94209 37820
rect 0 37568 80 37588
rect 0 37528 268 37568
rect 308 37528 317 37568
rect 0 37508 80 37528
rect 4343 37024 4352 37064
rect 4392 37024 4434 37064
rect 4474 37024 4516 37064
rect 4556 37024 4598 37064
rect 4638 37024 4680 37064
rect 4720 37024 4729 37064
rect 19463 37024 19472 37064
rect 19512 37024 19554 37064
rect 19594 37024 19636 37064
rect 19676 37024 19718 37064
rect 19758 37024 19800 37064
rect 19840 37024 19849 37064
rect 34583 37024 34592 37064
rect 34632 37024 34674 37064
rect 34714 37024 34756 37064
rect 34796 37024 34838 37064
rect 34878 37024 34920 37064
rect 34960 37024 34969 37064
rect 49703 37024 49712 37064
rect 49752 37024 49794 37064
rect 49834 37024 49876 37064
rect 49916 37024 49958 37064
rect 49998 37024 50040 37064
rect 50080 37024 50089 37064
rect 64823 37024 64832 37064
rect 64872 37024 64914 37064
rect 64954 37024 64996 37064
rect 65036 37024 65078 37064
rect 65118 37024 65160 37064
rect 65200 37024 65209 37064
rect 79943 37024 79952 37064
rect 79992 37024 80034 37064
rect 80074 37024 80116 37064
rect 80156 37024 80198 37064
rect 80238 37024 80280 37064
rect 80320 37024 80329 37064
rect 95063 37024 95072 37064
rect 95112 37024 95154 37064
rect 95194 37024 95236 37064
rect 95276 37024 95318 37064
rect 95358 37024 95400 37064
rect 95440 37024 95449 37064
rect 0 36728 80 36748
rect 0 36688 76 36728
rect 116 36688 125 36728
rect 0 36668 80 36688
rect 3103 36268 3112 36308
rect 3152 36268 3194 36308
rect 3234 36268 3276 36308
rect 3316 36268 3358 36308
rect 3398 36268 3440 36308
rect 3480 36268 3489 36308
rect 18223 36268 18232 36308
rect 18272 36268 18314 36308
rect 18354 36268 18396 36308
rect 18436 36268 18478 36308
rect 18518 36268 18560 36308
rect 18600 36268 18609 36308
rect 33343 36268 33352 36308
rect 33392 36268 33434 36308
rect 33474 36268 33516 36308
rect 33556 36268 33598 36308
rect 33638 36268 33680 36308
rect 33720 36268 33729 36308
rect 48463 36268 48472 36308
rect 48512 36268 48554 36308
rect 48594 36268 48636 36308
rect 48676 36268 48718 36308
rect 48758 36268 48800 36308
rect 48840 36268 48849 36308
rect 63583 36268 63592 36308
rect 63632 36268 63674 36308
rect 63714 36268 63756 36308
rect 63796 36268 63838 36308
rect 63878 36268 63920 36308
rect 63960 36268 63969 36308
rect 78703 36268 78712 36308
rect 78752 36268 78794 36308
rect 78834 36268 78876 36308
rect 78916 36268 78958 36308
rect 78998 36268 79040 36308
rect 79080 36268 79089 36308
rect 93823 36268 93832 36308
rect 93872 36268 93914 36308
rect 93954 36268 93996 36308
rect 94036 36268 94078 36308
rect 94118 36268 94160 36308
rect 94200 36268 94209 36308
rect 0 35828 80 35908
rect 4343 35512 4352 35552
rect 4392 35512 4434 35552
rect 4474 35512 4516 35552
rect 4556 35512 4598 35552
rect 4638 35512 4680 35552
rect 4720 35512 4729 35552
rect 19463 35512 19472 35552
rect 19512 35512 19554 35552
rect 19594 35512 19636 35552
rect 19676 35512 19718 35552
rect 19758 35512 19800 35552
rect 19840 35512 19849 35552
rect 34583 35512 34592 35552
rect 34632 35512 34674 35552
rect 34714 35512 34756 35552
rect 34796 35512 34838 35552
rect 34878 35512 34920 35552
rect 34960 35512 34969 35552
rect 49703 35512 49712 35552
rect 49752 35512 49794 35552
rect 49834 35512 49876 35552
rect 49916 35512 49958 35552
rect 49998 35512 50040 35552
rect 50080 35512 50089 35552
rect 64823 35512 64832 35552
rect 64872 35512 64914 35552
rect 64954 35512 64996 35552
rect 65036 35512 65078 35552
rect 65118 35512 65160 35552
rect 65200 35512 65209 35552
rect 79943 35512 79952 35552
rect 79992 35512 80034 35552
rect 80074 35512 80116 35552
rect 80156 35512 80198 35552
rect 80238 35512 80280 35552
rect 80320 35512 80329 35552
rect 95063 35512 95072 35552
rect 95112 35512 95154 35552
rect 95194 35512 95236 35552
rect 95276 35512 95318 35552
rect 95358 35512 95400 35552
rect 95440 35512 95449 35552
rect 835 35176 844 35216
rect 884 35176 23500 35216
rect 23540 35176 23549 35216
rect 0 35048 80 35068
rect 0 35008 652 35048
rect 692 35008 701 35048
rect 0 34988 80 35008
rect 3103 34756 3112 34796
rect 3152 34756 3194 34796
rect 3234 34756 3276 34796
rect 3316 34756 3358 34796
rect 3398 34756 3440 34796
rect 3480 34756 3489 34796
rect 18223 34756 18232 34796
rect 18272 34756 18314 34796
rect 18354 34756 18396 34796
rect 18436 34756 18478 34796
rect 18518 34756 18560 34796
rect 18600 34756 18609 34796
rect 33343 34756 33352 34796
rect 33392 34756 33434 34796
rect 33474 34756 33516 34796
rect 33556 34756 33598 34796
rect 33638 34756 33680 34796
rect 33720 34756 33729 34796
rect 48463 34756 48472 34796
rect 48512 34756 48554 34796
rect 48594 34756 48636 34796
rect 48676 34756 48718 34796
rect 48758 34756 48800 34796
rect 48840 34756 48849 34796
rect 63583 34756 63592 34796
rect 63632 34756 63674 34796
rect 63714 34756 63756 34796
rect 63796 34756 63838 34796
rect 63878 34756 63920 34796
rect 63960 34756 63969 34796
rect 78703 34756 78712 34796
rect 78752 34756 78794 34796
rect 78834 34756 78876 34796
rect 78916 34756 78958 34796
rect 78998 34756 79040 34796
rect 79080 34756 79089 34796
rect 93823 34756 93832 34796
rect 93872 34756 93914 34796
rect 93954 34756 93996 34796
rect 94036 34756 94078 34796
rect 94118 34756 94160 34796
rect 94200 34756 94209 34796
rect 835 34336 844 34376
rect 884 34336 29356 34376
rect 29396 34336 29405 34376
rect 0 34208 80 34228
rect 0 34168 652 34208
rect 692 34168 701 34208
rect 0 34148 80 34168
rect 4343 34000 4352 34040
rect 4392 34000 4434 34040
rect 4474 34000 4516 34040
rect 4556 34000 4598 34040
rect 4638 34000 4680 34040
rect 4720 34000 4729 34040
rect 19463 34000 19472 34040
rect 19512 34000 19554 34040
rect 19594 34000 19636 34040
rect 19676 34000 19718 34040
rect 19758 34000 19800 34040
rect 19840 34000 19849 34040
rect 34583 34000 34592 34040
rect 34632 34000 34674 34040
rect 34714 34000 34756 34040
rect 34796 34000 34838 34040
rect 34878 34000 34920 34040
rect 34960 34000 34969 34040
rect 49703 34000 49712 34040
rect 49752 34000 49794 34040
rect 49834 34000 49876 34040
rect 49916 34000 49958 34040
rect 49998 34000 50040 34040
rect 50080 34000 50089 34040
rect 64823 34000 64832 34040
rect 64872 34000 64914 34040
rect 64954 34000 64996 34040
rect 65036 34000 65078 34040
rect 65118 34000 65160 34040
rect 65200 34000 65209 34040
rect 79943 34000 79952 34040
rect 79992 34000 80034 34040
rect 80074 34000 80116 34040
rect 80156 34000 80198 34040
rect 80238 34000 80280 34040
rect 80320 34000 80329 34040
rect 95063 34000 95072 34040
rect 95112 34000 95154 34040
rect 95194 34000 95236 34040
rect 95276 34000 95318 34040
rect 95358 34000 95400 34040
rect 95440 34000 95449 34040
rect 835 33664 844 33704
rect 884 33664 29644 33704
rect 29684 33664 29693 33704
rect 0 33368 80 33388
rect 0 33328 652 33368
rect 692 33328 701 33368
rect 0 33308 80 33328
rect 3103 33244 3112 33284
rect 3152 33244 3194 33284
rect 3234 33244 3276 33284
rect 3316 33244 3358 33284
rect 3398 33244 3440 33284
rect 3480 33244 3489 33284
rect 18223 33244 18232 33284
rect 18272 33244 18314 33284
rect 18354 33244 18396 33284
rect 18436 33244 18478 33284
rect 18518 33244 18560 33284
rect 18600 33244 18609 33284
rect 33343 33244 33352 33284
rect 33392 33244 33434 33284
rect 33474 33244 33516 33284
rect 33556 33244 33598 33284
rect 33638 33244 33680 33284
rect 33720 33244 33729 33284
rect 48463 33244 48472 33284
rect 48512 33244 48554 33284
rect 48594 33244 48636 33284
rect 48676 33244 48718 33284
rect 48758 33244 48800 33284
rect 48840 33244 48849 33284
rect 63583 33244 63592 33284
rect 63632 33244 63674 33284
rect 63714 33244 63756 33284
rect 63796 33244 63838 33284
rect 63878 33244 63920 33284
rect 63960 33244 63969 33284
rect 78703 33244 78712 33284
rect 78752 33244 78794 33284
rect 78834 33244 78876 33284
rect 78916 33244 78958 33284
rect 78998 33244 79040 33284
rect 79080 33244 79089 33284
rect 93823 33244 93832 33284
rect 93872 33244 93914 33284
rect 93954 33244 93996 33284
rect 94036 33244 94078 33284
rect 94118 33244 94160 33284
rect 94200 33244 94209 33284
rect 835 32824 844 32864
rect 884 32824 29068 32864
rect 29108 32824 29117 32864
rect 0 32528 80 32548
rect 0 32488 652 32528
rect 692 32488 701 32528
rect 4343 32488 4352 32528
rect 4392 32488 4434 32528
rect 4474 32488 4516 32528
rect 4556 32488 4598 32528
rect 4638 32488 4680 32528
rect 4720 32488 4729 32528
rect 19463 32488 19472 32528
rect 19512 32488 19554 32528
rect 19594 32488 19636 32528
rect 19676 32488 19718 32528
rect 19758 32488 19800 32528
rect 19840 32488 19849 32528
rect 34583 32488 34592 32528
rect 34632 32488 34674 32528
rect 34714 32488 34756 32528
rect 34796 32488 34838 32528
rect 34878 32488 34920 32528
rect 34960 32488 34969 32528
rect 49703 32488 49712 32528
rect 49752 32488 49794 32528
rect 49834 32488 49876 32528
rect 49916 32488 49958 32528
rect 49998 32488 50040 32528
rect 50080 32488 50089 32528
rect 64823 32488 64832 32528
rect 64872 32488 64914 32528
rect 64954 32488 64996 32528
rect 65036 32488 65078 32528
rect 65118 32488 65160 32528
rect 65200 32488 65209 32528
rect 79943 32488 79952 32528
rect 79992 32488 80034 32528
rect 80074 32488 80116 32528
rect 80156 32488 80198 32528
rect 80238 32488 80280 32528
rect 80320 32488 80329 32528
rect 95063 32488 95072 32528
rect 95112 32488 95154 32528
rect 95194 32488 95236 32528
rect 95276 32488 95318 32528
rect 95358 32488 95400 32528
rect 95440 32488 95449 32528
rect 0 32468 80 32488
rect 27043 31900 27052 31940
rect 27092 31900 27532 31940
rect 27572 31900 27581 31940
rect 3103 31732 3112 31772
rect 3152 31732 3194 31772
rect 3234 31732 3276 31772
rect 3316 31732 3358 31772
rect 3398 31732 3440 31772
rect 3480 31732 3489 31772
rect 18223 31732 18232 31772
rect 18272 31732 18314 31772
rect 18354 31732 18396 31772
rect 18436 31732 18478 31772
rect 18518 31732 18560 31772
rect 18600 31732 18609 31772
rect 33343 31732 33352 31772
rect 33392 31732 33434 31772
rect 33474 31732 33516 31772
rect 33556 31732 33598 31772
rect 33638 31732 33680 31772
rect 33720 31732 33729 31772
rect 48463 31732 48472 31772
rect 48512 31732 48554 31772
rect 48594 31732 48636 31772
rect 48676 31732 48718 31772
rect 48758 31732 48800 31772
rect 48840 31732 48849 31772
rect 63583 31732 63592 31772
rect 63632 31732 63674 31772
rect 63714 31732 63756 31772
rect 63796 31732 63838 31772
rect 63878 31732 63920 31772
rect 63960 31732 63969 31772
rect 78703 31732 78712 31772
rect 78752 31732 78794 31772
rect 78834 31732 78876 31772
rect 78916 31732 78958 31772
rect 78998 31732 79040 31772
rect 79080 31732 79089 31772
rect 93823 31732 93832 31772
rect 93872 31732 93914 31772
rect 93954 31732 93996 31772
rect 94036 31732 94078 31772
rect 94118 31732 94160 31772
rect 94200 31732 94209 31772
rect 0 31688 80 31708
rect 0 31648 652 31688
rect 692 31648 701 31688
rect 0 31628 80 31648
rect 22627 31312 22636 31352
rect 22676 31312 27916 31352
rect 27956 31312 27965 31352
rect 21763 31228 21772 31268
rect 21812 31228 28780 31268
rect 28820 31228 28829 31268
rect 23779 31144 23788 31184
rect 23828 31144 27340 31184
rect 27380 31144 27389 31184
rect 4343 30976 4352 31016
rect 4392 30976 4434 31016
rect 4474 30976 4516 31016
rect 4556 30976 4598 31016
rect 4638 30976 4680 31016
rect 4720 30976 4729 31016
rect 19463 30976 19472 31016
rect 19512 30976 19554 31016
rect 19594 30976 19636 31016
rect 19676 30976 19718 31016
rect 19758 30976 19800 31016
rect 19840 30976 19849 31016
rect 34583 30976 34592 31016
rect 34632 30976 34674 31016
rect 34714 30976 34756 31016
rect 34796 30976 34838 31016
rect 34878 30976 34920 31016
rect 34960 30976 34969 31016
rect 49703 30976 49712 31016
rect 49752 30976 49794 31016
rect 49834 30976 49876 31016
rect 49916 30976 49958 31016
rect 49998 30976 50040 31016
rect 50080 30976 50089 31016
rect 64823 30976 64832 31016
rect 64872 30976 64914 31016
rect 64954 30976 64996 31016
rect 65036 30976 65078 31016
rect 65118 30976 65160 31016
rect 65200 30976 65209 31016
rect 79943 30976 79952 31016
rect 79992 30976 80034 31016
rect 80074 30976 80116 31016
rect 80156 30976 80198 31016
rect 80238 30976 80280 31016
rect 80320 30976 80329 31016
rect 95063 30976 95072 31016
rect 95112 30976 95154 31016
rect 95194 30976 95236 31016
rect 95276 30976 95318 31016
rect 95358 30976 95400 31016
rect 95440 30976 95449 31016
rect 0 30848 80 30868
rect 0 30808 652 30848
rect 692 30808 701 30848
rect 0 30788 80 30808
rect 26755 30640 26764 30680
rect 26804 30640 27628 30680
rect 27668 30640 27677 30680
rect 32803 30640 32812 30680
rect 32852 30640 33964 30680
rect 34004 30640 34013 30680
rect 28771 30556 28780 30596
rect 28820 30556 33100 30596
rect 33140 30556 34348 30596
rect 34388 30556 34397 30596
rect 35107 30388 35116 30428
rect 35156 30388 35596 30428
rect 35636 30388 35645 30428
rect 3103 30220 3112 30260
rect 3152 30220 3194 30260
rect 3234 30220 3276 30260
rect 3316 30220 3358 30260
rect 3398 30220 3440 30260
rect 3480 30220 3489 30260
rect 18223 30220 18232 30260
rect 18272 30220 18314 30260
rect 18354 30220 18396 30260
rect 18436 30220 18478 30260
rect 18518 30220 18560 30260
rect 18600 30220 18609 30260
rect 28291 30220 28300 30260
rect 28340 30220 29164 30260
rect 29204 30220 29213 30260
rect 31267 30220 31276 30260
rect 31316 30220 32716 30260
rect 32756 30220 32765 30260
rect 33343 30220 33352 30260
rect 33392 30220 33434 30260
rect 33474 30220 33516 30260
rect 33556 30220 33598 30260
rect 33638 30220 33680 30260
rect 33720 30220 33729 30260
rect 48463 30220 48472 30260
rect 48512 30220 48554 30260
rect 48594 30220 48636 30260
rect 48676 30220 48718 30260
rect 48758 30220 48800 30260
rect 48840 30220 48849 30260
rect 63583 30220 63592 30260
rect 63632 30220 63674 30260
rect 63714 30220 63756 30260
rect 63796 30220 63838 30260
rect 63878 30220 63920 30260
rect 63960 30220 63969 30260
rect 78703 30220 78712 30260
rect 78752 30220 78794 30260
rect 78834 30220 78876 30260
rect 78916 30220 78958 30260
rect 78998 30220 79040 30260
rect 79080 30220 79089 30260
rect 93823 30220 93832 30260
rect 93872 30220 93914 30260
rect 93954 30220 93996 30260
rect 94036 30220 94078 30260
rect 94118 30220 94160 30260
rect 94200 30220 94209 30260
rect 643 30052 652 30092
rect 692 30052 701 30092
rect 0 30008 80 30028
rect 652 30008 692 30052
rect 0 29968 692 30008
rect 0 29948 80 29968
rect 1123 29800 1132 29840
rect 1172 29800 19948 29840
rect 19988 29800 19997 29840
rect 4343 29464 4352 29504
rect 4392 29464 4434 29504
rect 4474 29464 4516 29504
rect 4556 29464 4598 29504
rect 4638 29464 4680 29504
rect 4720 29464 4729 29504
rect 19463 29464 19472 29504
rect 19512 29464 19554 29504
rect 19594 29464 19636 29504
rect 19676 29464 19718 29504
rect 19758 29464 19800 29504
rect 19840 29464 19849 29504
rect 34583 29464 34592 29504
rect 34632 29464 34674 29504
rect 34714 29464 34756 29504
rect 34796 29464 34838 29504
rect 34878 29464 34920 29504
rect 34960 29464 34969 29504
rect 49703 29464 49712 29504
rect 49752 29464 49794 29504
rect 49834 29464 49876 29504
rect 49916 29464 49958 29504
rect 49998 29464 50040 29504
rect 50080 29464 50089 29504
rect 64823 29464 64832 29504
rect 64872 29464 64914 29504
rect 64954 29464 64996 29504
rect 65036 29464 65078 29504
rect 65118 29464 65160 29504
rect 65200 29464 65209 29504
rect 79943 29464 79952 29504
rect 79992 29464 80034 29504
rect 80074 29464 80116 29504
rect 80156 29464 80198 29504
rect 80238 29464 80280 29504
rect 80320 29464 80329 29504
rect 95063 29464 95072 29504
rect 95112 29464 95154 29504
rect 95194 29464 95236 29504
rect 95276 29464 95318 29504
rect 95358 29464 95400 29504
rect 95440 29464 95449 29504
rect 0 29168 80 29188
rect 0 29128 652 29168
rect 692 29128 701 29168
rect 0 29108 80 29128
rect 35779 28960 35788 29000
rect 35828 28960 36460 29000
rect 36500 28960 36509 29000
rect 3103 28708 3112 28748
rect 3152 28708 3194 28748
rect 3234 28708 3276 28748
rect 3316 28708 3358 28748
rect 3398 28708 3440 28748
rect 3480 28708 3489 28748
rect 18223 28708 18232 28748
rect 18272 28708 18314 28748
rect 18354 28708 18396 28748
rect 18436 28708 18478 28748
rect 18518 28708 18560 28748
rect 18600 28708 18609 28748
rect 33343 28708 33352 28748
rect 33392 28708 33434 28748
rect 33474 28708 33516 28748
rect 33556 28708 33598 28748
rect 33638 28708 33680 28748
rect 33720 28708 33729 28748
rect 48463 28708 48472 28748
rect 48512 28708 48554 28748
rect 48594 28708 48636 28748
rect 48676 28708 48718 28748
rect 48758 28708 48800 28748
rect 48840 28708 48849 28748
rect 63583 28708 63592 28748
rect 63632 28708 63674 28748
rect 63714 28708 63756 28748
rect 63796 28708 63838 28748
rect 63878 28708 63920 28748
rect 63960 28708 63969 28748
rect 78703 28708 78712 28748
rect 78752 28708 78794 28748
rect 78834 28708 78876 28748
rect 78916 28708 78958 28748
rect 78998 28708 79040 28748
rect 79080 28708 79089 28748
rect 93823 28708 93832 28748
rect 93872 28708 93914 28748
rect 93954 28708 93996 28748
rect 94036 28708 94078 28748
rect 94118 28708 94160 28748
rect 94200 28708 94209 28748
rect 21379 28540 21388 28580
rect 21428 28540 22060 28580
rect 22100 28540 22109 28580
rect 28195 28456 28204 28496
rect 28244 28456 28780 28496
rect 28820 28456 28829 28496
rect 23920 28372 27532 28412
rect 27572 28372 27581 28412
rect 0 28328 80 28348
rect 23920 28328 23960 28372
rect 0 28288 652 28328
rect 692 28288 701 28328
rect 835 28288 844 28328
rect 884 28288 6320 28328
rect 15331 28288 15340 28328
rect 15380 28288 22444 28328
rect 22484 28288 23212 28328
rect 23252 28288 23261 28328
rect 23395 28288 23404 28328
rect 23444 28288 23960 28328
rect 27139 28288 27148 28328
rect 27188 28288 28108 28328
rect 28148 28288 31180 28328
rect 31220 28288 31229 28328
rect 0 28268 80 28288
rect 6280 28244 6320 28288
rect 6280 28204 28012 28244
rect 28052 28204 28061 28244
rect 23491 28120 23500 28160
rect 23540 28120 26860 28160
rect 26900 28120 26909 28160
rect 28483 28120 28492 28160
rect 28532 28120 29452 28160
rect 29492 28120 29501 28160
rect 18211 28036 18220 28076
rect 18260 28036 23404 28076
rect 23444 28036 23453 28076
rect 4343 27952 4352 27992
rect 4392 27952 4434 27992
rect 4474 27952 4516 27992
rect 4556 27952 4598 27992
rect 4638 27952 4680 27992
rect 4720 27952 4729 27992
rect 19463 27952 19472 27992
rect 19512 27952 19554 27992
rect 19594 27952 19636 27992
rect 19676 27952 19718 27992
rect 19758 27952 19800 27992
rect 19840 27952 19849 27992
rect 34583 27952 34592 27992
rect 34632 27952 34674 27992
rect 34714 27952 34756 27992
rect 34796 27952 34838 27992
rect 34878 27952 34920 27992
rect 34960 27952 34969 27992
rect 49703 27952 49712 27992
rect 49752 27952 49794 27992
rect 49834 27952 49876 27992
rect 49916 27952 49958 27992
rect 49998 27952 50040 27992
rect 50080 27952 50089 27992
rect 64823 27952 64832 27992
rect 64872 27952 64914 27992
rect 64954 27952 64996 27992
rect 65036 27952 65078 27992
rect 65118 27952 65160 27992
rect 65200 27952 65209 27992
rect 79943 27952 79952 27992
rect 79992 27952 80034 27992
rect 80074 27952 80116 27992
rect 80156 27952 80198 27992
rect 80238 27952 80280 27992
rect 80320 27952 80329 27992
rect 95063 27952 95072 27992
rect 95112 27952 95154 27992
rect 95194 27952 95236 27992
rect 95276 27952 95318 27992
rect 95358 27952 95400 27992
rect 95440 27952 95449 27992
rect 739 27784 748 27824
rect 788 27784 20044 27824
rect 20084 27784 21484 27824
rect 21524 27784 21533 27824
rect 22339 27784 22348 27824
rect 22388 27784 23308 27824
rect 23348 27784 28300 27824
rect 28340 27784 28349 27824
rect 21571 27700 21580 27740
rect 21620 27700 22540 27740
rect 22580 27700 23404 27740
rect 23444 27700 23453 27740
rect 26563 27700 26572 27740
rect 26612 27700 28396 27740
rect 28436 27700 28445 27740
rect 29443 27700 29452 27740
rect 29492 27700 29684 27740
rect 29644 27656 29684 27700
rect 17251 27616 17260 27656
rect 17300 27616 18124 27656
rect 18164 27616 18173 27656
rect 18499 27616 18508 27656
rect 18548 27616 20236 27656
rect 20276 27616 20285 27656
rect 26371 27616 26380 27656
rect 26420 27616 26956 27656
rect 26996 27616 27005 27656
rect 29635 27616 29644 27656
rect 29684 27616 29693 27656
rect 29155 27532 29164 27572
rect 29204 27532 29452 27572
rect 29492 27532 30028 27572
rect 30068 27532 30077 27572
rect 0 27488 80 27508
rect 0 27448 652 27488
rect 692 27448 701 27488
rect 931 27448 940 27488
rect 980 27448 20140 27488
rect 20180 27448 21676 27488
rect 21716 27448 21725 27488
rect 28099 27448 28108 27488
rect 28148 27448 29260 27488
rect 29300 27448 29309 27488
rect 0 27428 80 27448
rect 23587 27364 23596 27404
rect 23636 27364 23960 27404
rect 29347 27364 29356 27404
rect 29396 27364 30124 27404
rect 30164 27364 30173 27404
rect 23920 27320 23960 27364
rect 23920 27280 34924 27320
rect 34964 27280 34973 27320
rect 3103 27196 3112 27236
rect 3152 27196 3194 27236
rect 3234 27196 3276 27236
rect 3316 27196 3358 27236
rect 3398 27196 3440 27236
rect 3480 27196 3489 27236
rect 18223 27196 18232 27236
rect 18272 27196 18314 27236
rect 18354 27196 18396 27236
rect 18436 27196 18478 27236
rect 18518 27196 18560 27236
rect 18600 27196 18609 27236
rect 33343 27196 33352 27236
rect 33392 27196 33434 27236
rect 33474 27196 33516 27236
rect 33556 27196 33598 27236
rect 33638 27196 33680 27236
rect 33720 27196 33729 27236
rect 48463 27196 48472 27236
rect 48512 27196 48554 27236
rect 48594 27196 48636 27236
rect 48676 27196 48718 27236
rect 48758 27196 48800 27236
rect 48840 27196 48849 27236
rect 63583 27196 63592 27236
rect 63632 27196 63674 27236
rect 63714 27196 63756 27236
rect 63796 27196 63838 27236
rect 63878 27196 63920 27236
rect 63960 27196 63969 27236
rect 78703 27196 78712 27236
rect 78752 27196 78794 27236
rect 78834 27196 78876 27236
rect 78916 27196 78958 27236
rect 78998 27196 79040 27236
rect 79080 27196 79089 27236
rect 93823 27196 93832 27236
rect 93872 27196 93914 27236
rect 93954 27196 93996 27236
rect 94036 27196 94078 27236
rect 94118 27196 94160 27236
rect 94200 27196 94209 27236
rect 35875 27028 35884 27068
rect 35924 27028 37324 27068
rect 37364 27028 37373 27068
rect 1027 26944 1036 26984
rect 1076 26944 19948 26984
rect 19988 26944 19997 26984
rect 20227 26860 20236 26900
rect 20276 26860 20428 26900
rect 20468 26860 25804 26900
rect 25844 26860 26380 26900
rect 26420 26860 26429 26900
rect 20131 26776 20140 26816
rect 20180 26776 20620 26816
rect 20660 26776 21772 26816
rect 21812 26776 21821 26816
rect 35395 26776 35404 26816
rect 35444 26776 36172 26816
rect 36212 26776 36221 26816
rect 0 26648 80 26668
rect 0 26608 652 26648
rect 692 26608 701 26648
rect 14851 26608 14860 26648
rect 14900 26608 20332 26648
rect 20372 26608 20381 26648
rect 0 26588 80 26608
rect 4343 26440 4352 26480
rect 4392 26440 4434 26480
rect 4474 26440 4516 26480
rect 4556 26440 4598 26480
rect 4638 26440 4680 26480
rect 4720 26440 4729 26480
rect 19463 26440 19472 26480
rect 19512 26440 19554 26480
rect 19594 26440 19636 26480
rect 19676 26440 19718 26480
rect 19758 26440 19800 26480
rect 19840 26440 19849 26480
rect 34583 26440 34592 26480
rect 34632 26440 34674 26480
rect 34714 26440 34756 26480
rect 34796 26440 34838 26480
rect 34878 26440 34920 26480
rect 34960 26440 34969 26480
rect 49703 26440 49712 26480
rect 49752 26440 49794 26480
rect 49834 26440 49876 26480
rect 49916 26440 49958 26480
rect 49998 26440 50040 26480
rect 50080 26440 50089 26480
rect 64823 26440 64832 26480
rect 64872 26440 64914 26480
rect 64954 26440 64996 26480
rect 65036 26440 65078 26480
rect 65118 26440 65160 26480
rect 65200 26440 65209 26480
rect 79943 26440 79952 26480
rect 79992 26440 80034 26480
rect 80074 26440 80116 26480
rect 80156 26440 80198 26480
rect 80238 26440 80280 26480
rect 80320 26440 80329 26480
rect 95063 26440 95072 26480
rect 95112 26440 95154 26480
rect 95194 26440 95236 26480
rect 95276 26440 95318 26480
rect 95358 26440 95400 26480
rect 95440 26440 95449 26480
rect 16099 26356 16108 26396
rect 16148 26356 16588 26396
rect 16628 26356 22636 26396
rect 22676 26356 22685 26396
rect 259 26188 268 26228
rect 308 26188 23960 26228
rect 23920 26144 23960 26188
rect 23920 26104 39628 26144
rect 39668 26104 39677 26144
rect 25987 26020 25996 26060
rect 26036 26020 26380 26060
rect 26420 26020 26429 26060
rect 26851 26020 26860 26060
rect 26900 26020 28204 26060
rect 28244 26020 28253 26060
rect 35299 26020 35308 26060
rect 35348 26020 35500 26060
rect 35540 26020 35549 26060
rect 0 25808 80 25828
rect 0 25768 652 25808
rect 692 25768 701 25808
rect 0 25748 80 25768
rect 3103 25684 3112 25724
rect 3152 25684 3194 25724
rect 3234 25684 3276 25724
rect 3316 25684 3358 25724
rect 3398 25684 3440 25724
rect 3480 25684 3489 25724
rect 18223 25684 18232 25724
rect 18272 25684 18314 25724
rect 18354 25684 18396 25724
rect 18436 25684 18478 25724
rect 18518 25684 18560 25724
rect 18600 25684 18609 25724
rect 33343 25684 33352 25724
rect 33392 25684 33434 25724
rect 33474 25684 33516 25724
rect 33556 25684 33598 25724
rect 33638 25684 33680 25724
rect 33720 25684 33729 25724
rect 48463 25684 48472 25724
rect 48512 25684 48554 25724
rect 48594 25684 48636 25724
rect 48676 25684 48718 25724
rect 48758 25684 48800 25724
rect 48840 25684 48849 25724
rect 63583 25684 63592 25724
rect 63632 25684 63674 25724
rect 63714 25684 63756 25724
rect 63796 25684 63838 25724
rect 63878 25684 63920 25724
rect 63960 25684 63969 25724
rect 78703 25684 78712 25724
rect 78752 25684 78794 25724
rect 78834 25684 78876 25724
rect 78916 25684 78958 25724
rect 78998 25684 79040 25724
rect 79080 25684 79089 25724
rect 93823 25684 93832 25724
rect 93872 25684 93914 25724
rect 93954 25684 93996 25724
rect 94036 25684 94078 25724
rect 94118 25684 94160 25724
rect 94200 25684 94209 25724
rect 26371 25516 26380 25556
rect 26420 25516 28204 25556
rect 28244 25516 28253 25556
rect 931 25432 940 25472
rect 980 25432 6320 25472
rect 6280 25304 6320 25432
rect 6280 25264 28396 25304
rect 28436 25264 29260 25304
rect 29300 25264 30028 25304
rect 30068 25264 30077 25304
rect 35203 25180 35212 25220
rect 35252 25180 35596 25220
rect 35636 25180 35645 25220
rect 28003 25096 28012 25136
rect 28052 25096 28492 25136
rect 28532 25096 28541 25136
rect 0 24968 80 24988
rect 0 24928 652 24968
rect 692 24928 701 24968
rect 4343 24928 4352 24968
rect 4392 24928 4434 24968
rect 4474 24928 4516 24968
rect 4556 24928 4598 24968
rect 4638 24928 4680 24968
rect 4720 24928 4729 24968
rect 19463 24928 19472 24968
rect 19512 24928 19554 24968
rect 19594 24928 19636 24968
rect 19676 24928 19718 24968
rect 19758 24928 19800 24968
rect 19840 24928 19849 24968
rect 34583 24928 34592 24968
rect 34632 24928 34674 24968
rect 34714 24928 34756 24968
rect 34796 24928 34838 24968
rect 34878 24928 34920 24968
rect 34960 24928 34969 24968
rect 49703 24928 49712 24968
rect 49752 24928 49794 24968
rect 49834 24928 49876 24968
rect 49916 24928 49958 24968
rect 49998 24928 50040 24968
rect 50080 24928 50089 24968
rect 64823 24928 64832 24968
rect 64872 24928 64914 24968
rect 64954 24928 64996 24968
rect 65036 24928 65078 24968
rect 65118 24928 65160 24968
rect 65200 24928 65209 24968
rect 79943 24928 79952 24968
rect 79992 24928 80034 24968
rect 80074 24928 80116 24968
rect 80156 24928 80198 24968
rect 80238 24928 80280 24968
rect 80320 24928 80329 24968
rect 95063 24928 95072 24968
rect 95112 24928 95154 24968
rect 95194 24928 95236 24968
rect 95276 24928 95318 24968
rect 95358 24928 95400 24968
rect 95440 24928 95449 24968
rect 0 24908 80 24928
rect 22627 24592 22636 24632
rect 22676 24592 23020 24632
rect 23060 24592 23069 24632
rect 27523 24508 27532 24548
rect 27572 24508 29836 24548
rect 29876 24508 35212 24548
rect 35252 24508 35261 24548
rect 3103 24172 3112 24212
rect 3152 24172 3194 24212
rect 3234 24172 3276 24212
rect 3316 24172 3358 24212
rect 3398 24172 3440 24212
rect 3480 24172 3489 24212
rect 18223 24172 18232 24212
rect 18272 24172 18314 24212
rect 18354 24172 18396 24212
rect 18436 24172 18478 24212
rect 18518 24172 18560 24212
rect 18600 24172 18609 24212
rect 33343 24172 33352 24212
rect 33392 24172 33434 24212
rect 33474 24172 33516 24212
rect 33556 24172 33598 24212
rect 33638 24172 33680 24212
rect 33720 24172 33729 24212
rect 48463 24172 48472 24212
rect 48512 24172 48554 24212
rect 48594 24172 48636 24212
rect 48676 24172 48718 24212
rect 48758 24172 48800 24212
rect 48840 24172 48849 24212
rect 63583 24172 63592 24212
rect 63632 24172 63674 24212
rect 63714 24172 63756 24212
rect 63796 24172 63838 24212
rect 63878 24172 63920 24212
rect 63960 24172 63969 24212
rect 78703 24172 78712 24212
rect 78752 24172 78794 24212
rect 78834 24172 78876 24212
rect 78916 24172 78958 24212
rect 78998 24172 79040 24212
rect 79080 24172 79089 24212
rect 93823 24172 93832 24212
rect 93872 24172 93914 24212
rect 93954 24172 93996 24212
rect 94036 24172 94078 24212
rect 94118 24172 94160 24212
rect 94200 24172 94209 24212
rect 0 24128 80 24148
rect 0 24088 652 24128
rect 692 24088 701 24128
rect 0 24068 80 24088
rect 25411 23836 25420 23876
rect 25460 23836 32812 23876
rect 32852 23836 32861 23876
rect 35491 23836 35500 23876
rect 35540 23836 39916 23876
rect 39956 23836 39965 23876
rect 35500 23792 35540 23836
rect 835 23752 844 23792
rect 884 23752 30124 23792
rect 30164 23752 30173 23792
rect 34435 23752 34444 23792
rect 34484 23752 35540 23792
rect 28483 23668 28492 23708
rect 28532 23668 28972 23708
rect 29012 23668 29644 23708
rect 29684 23668 29693 23708
rect 32803 23584 32812 23624
rect 32852 23584 33772 23624
rect 33812 23584 35404 23624
rect 35444 23584 35453 23624
rect 4343 23416 4352 23456
rect 4392 23416 4434 23456
rect 4474 23416 4516 23456
rect 4556 23416 4598 23456
rect 4638 23416 4680 23456
rect 4720 23416 4729 23456
rect 19463 23416 19472 23456
rect 19512 23416 19554 23456
rect 19594 23416 19636 23456
rect 19676 23416 19718 23456
rect 19758 23416 19800 23456
rect 19840 23416 19849 23456
rect 34583 23416 34592 23456
rect 34632 23416 34674 23456
rect 34714 23416 34756 23456
rect 34796 23416 34838 23456
rect 34878 23416 34920 23456
rect 34960 23416 34969 23456
rect 49703 23416 49712 23456
rect 49752 23416 49794 23456
rect 49834 23416 49876 23456
rect 49916 23416 49958 23456
rect 49998 23416 50040 23456
rect 50080 23416 50089 23456
rect 64823 23416 64832 23456
rect 64872 23416 64914 23456
rect 64954 23416 64996 23456
rect 65036 23416 65078 23456
rect 65118 23416 65160 23456
rect 65200 23416 65209 23456
rect 79943 23416 79952 23456
rect 79992 23416 80034 23456
rect 80074 23416 80116 23456
rect 80156 23416 80198 23456
rect 80238 23416 80280 23456
rect 80320 23416 80329 23456
rect 95063 23416 95072 23456
rect 95112 23416 95154 23456
rect 95194 23416 95236 23456
rect 95276 23416 95318 23456
rect 95358 23416 95400 23456
rect 95440 23416 95449 23456
rect 0 23288 80 23308
rect 0 23248 652 23288
rect 692 23248 701 23288
rect 0 23228 80 23248
rect 15235 23080 15244 23120
rect 15284 23080 19756 23120
rect 19796 23080 21868 23120
rect 21908 23080 24556 23120
rect 24596 23080 24605 23120
rect 35299 23080 35308 23120
rect 35348 23080 40396 23120
rect 40436 23080 40445 23120
rect 21763 22828 21772 22868
rect 21812 22828 28588 22868
rect 28628 22828 28637 22868
rect 3103 22660 3112 22700
rect 3152 22660 3194 22700
rect 3234 22660 3276 22700
rect 3316 22660 3358 22700
rect 3398 22660 3440 22700
rect 3480 22660 3489 22700
rect 18223 22660 18232 22700
rect 18272 22660 18314 22700
rect 18354 22660 18396 22700
rect 18436 22660 18478 22700
rect 18518 22660 18560 22700
rect 18600 22660 18609 22700
rect 33343 22660 33352 22700
rect 33392 22660 33434 22700
rect 33474 22660 33516 22700
rect 33556 22660 33598 22700
rect 33638 22660 33680 22700
rect 33720 22660 33729 22700
rect 39523 22660 39532 22700
rect 39572 22660 39916 22700
rect 39956 22660 39965 22700
rect 48463 22660 48472 22700
rect 48512 22660 48554 22700
rect 48594 22660 48636 22700
rect 48676 22660 48718 22700
rect 48758 22660 48800 22700
rect 48840 22660 48849 22700
rect 63583 22660 63592 22700
rect 63632 22660 63674 22700
rect 63714 22660 63756 22700
rect 63796 22660 63838 22700
rect 63878 22660 63920 22700
rect 63960 22660 63969 22700
rect 78703 22660 78712 22700
rect 78752 22660 78794 22700
rect 78834 22660 78876 22700
rect 78916 22660 78958 22700
rect 78998 22660 79040 22700
rect 79080 22660 79089 22700
rect 93823 22660 93832 22700
rect 93872 22660 93914 22700
rect 93954 22660 93996 22700
rect 94036 22660 94078 22700
rect 94118 22660 94160 22700
rect 94200 22660 94209 22700
rect 28867 22576 28876 22616
rect 28916 22576 34156 22616
rect 34196 22576 34924 22616
rect 34964 22576 34973 22616
rect 27235 22492 27244 22532
rect 27284 22492 32620 22532
rect 32660 22492 32780 22532
rect 0 22388 80 22468
rect 32740 22448 32780 22492
rect 28675 22408 28684 22448
rect 28724 22408 28876 22448
rect 28916 22408 29164 22448
rect 29204 22408 29213 22448
rect 32740 22408 35596 22448
rect 35636 22408 35980 22448
rect 36020 22408 36029 22448
rect 26563 22324 26572 22364
rect 26612 22324 28780 22364
rect 28820 22324 28829 22364
rect 32515 22240 32524 22280
rect 32564 22240 34060 22280
rect 34100 22240 34109 22280
rect 23395 22156 23404 22196
rect 23444 22156 24172 22196
rect 24212 22156 24221 22196
rect 34156 22112 34196 22408
rect 34339 22324 34348 22364
rect 34388 22324 34732 22364
rect 34772 22324 35308 22364
rect 35348 22324 35357 22364
rect 35779 22324 35788 22364
rect 35828 22324 41548 22364
rect 41588 22324 41597 22364
rect 35395 22240 35404 22280
rect 35444 22240 36460 22280
rect 36500 22240 36509 22280
rect 34243 22156 34252 22196
rect 34292 22156 34868 22196
rect 35011 22156 35020 22196
rect 35060 22156 35692 22196
rect 35732 22156 35741 22196
rect 34828 22112 34868 22156
rect 17347 22072 17356 22112
rect 17396 22072 32428 22112
rect 32468 22072 32477 22112
rect 34147 22072 34156 22112
rect 34196 22072 34205 22112
rect 34348 22072 34636 22112
rect 34676 22072 34685 22112
rect 34819 22072 34828 22112
rect 34868 22072 34877 22112
rect 34348 21944 34388 22072
rect 34828 22028 34868 22072
rect 34828 21988 35020 22028
rect 35060 21988 35069 22028
rect 4343 21904 4352 21944
rect 4392 21904 4434 21944
rect 4474 21904 4516 21944
rect 4556 21904 4598 21944
rect 4638 21904 4680 21944
rect 4720 21904 4729 21944
rect 19463 21904 19472 21944
rect 19512 21904 19554 21944
rect 19594 21904 19636 21944
rect 19676 21904 19718 21944
rect 19758 21904 19800 21944
rect 19840 21904 19849 21944
rect 34339 21904 34348 21944
rect 34388 21904 34397 21944
rect 34583 21904 34592 21944
rect 34632 21904 34674 21944
rect 34714 21904 34756 21944
rect 34796 21904 34838 21944
rect 34878 21904 34920 21944
rect 34960 21904 34969 21944
rect 49703 21904 49712 21944
rect 49752 21904 49794 21944
rect 49834 21904 49876 21944
rect 49916 21904 49958 21944
rect 49998 21904 50040 21944
rect 50080 21904 50089 21944
rect 64823 21904 64832 21944
rect 64872 21904 64914 21944
rect 64954 21904 64996 21944
rect 65036 21904 65078 21944
rect 65118 21904 65160 21944
rect 65200 21904 65209 21944
rect 79943 21904 79952 21944
rect 79992 21904 80034 21944
rect 80074 21904 80116 21944
rect 80156 21904 80198 21944
rect 80238 21904 80280 21944
rect 80320 21904 80329 21944
rect 95063 21904 95072 21944
rect 95112 21904 95154 21944
rect 95194 21904 95236 21944
rect 95276 21904 95318 21944
rect 95358 21904 95400 21944
rect 95440 21904 95449 21944
rect 33091 21820 33100 21860
rect 33140 21820 35212 21860
rect 35252 21820 35261 21860
rect 76 21652 652 21692
rect 692 21652 701 21692
rect 76 21628 116 21652
rect 0 21568 116 21628
rect 163 21568 172 21608
rect 212 21568 28396 21608
rect 28436 21568 28445 21608
rect 29347 21568 29356 21608
rect 29396 21568 33196 21608
rect 33236 21568 33245 21608
rect 0 21548 80 21568
rect 29356 21524 29396 21568
rect 23971 21484 23980 21524
rect 24020 21484 24172 21524
rect 24212 21484 29396 21524
rect 3103 21148 3112 21188
rect 3152 21148 3194 21188
rect 3234 21148 3276 21188
rect 3316 21148 3358 21188
rect 3398 21148 3440 21188
rect 3480 21148 3489 21188
rect 18223 21148 18232 21188
rect 18272 21148 18314 21188
rect 18354 21148 18396 21188
rect 18436 21148 18478 21188
rect 18518 21148 18560 21188
rect 18600 21148 18609 21188
rect 33343 21148 33352 21188
rect 33392 21148 33434 21188
rect 33474 21148 33516 21188
rect 33556 21148 33598 21188
rect 33638 21148 33680 21188
rect 33720 21148 33729 21188
rect 48463 21148 48472 21188
rect 48512 21148 48554 21188
rect 48594 21148 48636 21188
rect 48676 21148 48718 21188
rect 48758 21148 48800 21188
rect 48840 21148 48849 21188
rect 63583 21148 63592 21188
rect 63632 21148 63674 21188
rect 63714 21148 63756 21188
rect 63796 21148 63838 21188
rect 63878 21148 63920 21188
rect 63960 21148 63969 21188
rect 78703 21148 78712 21188
rect 78752 21148 78794 21188
rect 78834 21148 78876 21188
rect 78916 21148 78958 21188
rect 78998 21148 79040 21188
rect 79080 21148 79089 21188
rect 93823 21148 93832 21188
rect 93872 21148 93914 21188
rect 93954 21148 93996 21188
rect 94036 21148 94078 21188
rect 94118 21148 94160 21188
rect 94200 21148 94209 21188
rect 29155 20896 29164 20936
rect 29204 20896 30316 20936
rect 30356 20896 30365 20936
rect 28867 20812 28876 20852
rect 28916 20812 31372 20852
rect 31412 20812 31421 20852
rect 0 20768 80 20788
rect 0 20728 652 20768
rect 692 20728 701 20768
rect 931 20728 940 20768
rect 980 20728 17740 20768
rect 17780 20728 19564 20768
rect 19604 20728 20140 20768
rect 20180 20728 20189 20768
rect 22627 20728 22636 20768
rect 22676 20728 23212 20768
rect 23252 20728 23261 20768
rect 29251 20728 29260 20768
rect 29300 20728 29644 20768
rect 29684 20728 30508 20768
rect 30548 20728 30557 20768
rect 0 20708 80 20728
rect 22915 20644 22924 20684
rect 22964 20644 34060 20684
rect 34100 20644 34109 20684
rect 23920 20560 30892 20600
rect 30932 20560 30941 20600
rect 23920 20516 23960 20560
rect 1123 20476 1132 20516
rect 1172 20476 23960 20516
rect 4343 20392 4352 20432
rect 4392 20392 4434 20432
rect 4474 20392 4516 20432
rect 4556 20392 4598 20432
rect 4638 20392 4680 20432
rect 4720 20392 4729 20432
rect 19463 20392 19472 20432
rect 19512 20392 19554 20432
rect 19594 20392 19636 20432
rect 19676 20392 19718 20432
rect 19758 20392 19800 20432
rect 19840 20392 19849 20432
rect 34583 20392 34592 20432
rect 34632 20392 34674 20432
rect 34714 20392 34756 20432
rect 34796 20392 34838 20432
rect 34878 20392 34920 20432
rect 34960 20392 34969 20432
rect 49703 20392 49712 20432
rect 49752 20392 49794 20432
rect 49834 20392 49876 20432
rect 49916 20392 49958 20432
rect 49998 20392 50040 20432
rect 50080 20392 50089 20432
rect 64823 20392 64832 20432
rect 64872 20392 64914 20432
rect 64954 20392 64996 20432
rect 65036 20392 65078 20432
rect 65118 20392 65160 20432
rect 65200 20392 65209 20432
rect 79943 20392 79952 20432
rect 79992 20392 80034 20432
rect 80074 20392 80116 20432
rect 80156 20392 80198 20432
rect 80238 20392 80280 20432
rect 80320 20392 80329 20432
rect 95063 20392 95072 20432
rect 95112 20392 95154 20432
rect 95194 20392 95236 20432
rect 95276 20392 95318 20432
rect 95358 20392 95400 20432
rect 95440 20392 95449 20432
rect 22051 20308 22060 20348
rect 22100 20308 22732 20348
rect 22772 20308 22781 20348
rect 23107 20224 23116 20264
rect 23156 20224 23165 20264
rect 23116 20180 23156 20224
rect 14947 20140 14956 20180
rect 14996 20140 15436 20180
rect 15476 20140 15485 20180
rect 20131 20140 20140 20180
rect 20180 20140 21772 20180
rect 21812 20140 22348 20180
rect 22388 20140 23500 20180
rect 23540 20140 23549 20180
rect 28099 20140 28108 20180
rect 28148 20140 29452 20180
rect 29492 20140 33812 20180
rect 33772 20096 33812 20140
rect 19459 20056 19468 20096
rect 19508 20056 21388 20096
rect 21428 20056 21868 20096
rect 21908 20056 21917 20096
rect 33763 20056 33772 20096
rect 33812 20056 34828 20096
rect 34868 20056 34877 20096
rect 35011 20056 35020 20096
rect 35060 20056 39916 20096
rect 39956 20056 41164 20096
rect 41204 20056 41213 20096
rect 739 19972 748 20012
rect 788 19972 15916 20012
rect 15956 19972 15965 20012
rect 0 19928 80 19948
rect 0 19888 652 19928
rect 692 19888 701 19928
rect 6280 19888 15628 19928
rect 15668 19888 15677 19928
rect 21379 19888 21388 19928
rect 21428 19888 22732 19928
rect 22772 19888 23308 19928
rect 23348 19888 23357 19928
rect 0 19868 80 19888
rect 6280 19844 6320 19888
rect 547 19804 556 19844
rect 596 19804 6320 19844
rect 37219 19804 37228 19844
rect 37268 19804 39244 19844
rect 39284 19804 39293 19844
rect 3103 19636 3112 19676
rect 3152 19636 3194 19676
rect 3234 19636 3276 19676
rect 3316 19636 3358 19676
rect 3398 19636 3440 19676
rect 3480 19636 3489 19676
rect 18223 19636 18232 19676
rect 18272 19636 18314 19676
rect 18354 19636 18396 19676
rect 18436 19636 18478 19676
rect 18518 19636 18560 19676
rect 18600 19636 18609 19676
rect 33343 19636 33352 19676
rect 33392 19636 33434 19676
rect 33474 19636 33516 19676
rect 33556 19636 33598 19676
rect 33638 19636 33680 19676
rect 33720 19636 33729 19676
rect 48463 19636 48472 19676
rect 48512 19636 48554 19676
rect 48594 19636 48636 19676
rect 48676 19636 48718 19676
rect 48758 19636 48800 19676
rect 48840 19636 48849 19676
rect 63583 19636 63592 19676
rect 63632 19636 63674 19676
rect 63714 19636 63756 19676
rect 63796 19636 63838 19676
rect 63878 19636 63920 19676
rect 63960 19636 63969 19676
rect 78703 19636 78712 19676
rect 78752 19636 78794 19676
rect 78834 19636 78876 19676
rect 78916 19636 78958 19676
rect 78998 19636 79040 19676
rect 79080 19636 79089 19676
rect 93823 19636 93832 19676
rect 93872 19636 93914 19676
rect 93954 19636 93996 19676
rect 94036 19636 94078 19676
rect 94118 19636 94160 19676
rect 94200 19636 94209 19676
rect 1027 19468 1036 19508
rect 1076 19468 18028 19508
rect 18068 19468 19468 19508
rect 19508 19468 19517 19508
rect 37507 19384 37516 19424
rect 37556 19384 38764 19424
rect 38804 19384 38813 19424
rect 19171 19300 19180 19340
rect 19220 19300 19372 19340
rect 19412 19300 21100 19340
rect 21140 19300 21149 19340
rect 23920 19300 37036 19340
rect 37076 19300 37085 19340
rect 23920 19256 23960 19300
rect 15907 19216 15916 19256
rect 15956 19216 16108 19256
rect 16148 19216 19660 19256
rect 19700 19216 21292 19256
rect 21332 19216 21341 19256
rect 23491 19216 23500 19256
rect 23540 19216 23960 19256
rect 33859 19216 33868 19256
rect 33908 19216 38860 19256
rect 38900 19216 40012 19256
rect 40052 19216 40061 19256
rect 15715 19132 15724 19172
rect 15764 19132 19084 19172
rect 19124 19132 22540 19172
rect 22580 19132 22589 19172
rect 0 19088 80 19108
rect 0 19048 652 19088
rect 692 19048 701 19088
rect 38755 19048 38764 19088
rect 38804 19048 39148 19088
rect 39188 19048 39532 19088
rect 39572 19048 39581 19088
rect 0 19028 80 19048
rect 4343 18880 4352 18920
rect 4392 18880 4434 18920
rect 4474 18880 4516 18920
rect 4556 18880 4598 18920
rect 4638 18880 4680 18920
rect 4720 18880 4729 18920
rect 19463 18880 19472 18920
rect 19512 18880 19554 18920
rect 19594 18880 19636 18920
rect 19676 18880 19718 18920
rect 19758 18880 19800 18920
rect 19840 18880 19849 18920
rect 32611 18880 32620 18920
rect 32660 18880 33868 18920
rect 33908 18880 33917 18920
rect 34583 18880 34592 18920
rect 34632 18880 34674 18920
rect 34714 18880 34756 18920
rect 34796 18880 34838 18920
rect 34878 18880 34920 18920
rect 34960 18880 34969 18920
rect 49703 18880 49712 18920
rect 49752 18880 49794 18920
rect 49834 18880 49876 18920
rect 49916 18880 49958 18920
rect 49998 18880 50040 18920
rect 50080 18880 50089 18920
rect 64823 18880 64832 18920
rect 64872 18880 64914 18920
rect 64954 18880 64996 18920
rect 65036 18880 65078 18920
rect 65118 18880 65160 18920
rect 65200 18880 65209 18920
rect 79943 18880 79952 18920
rect 79992 18880 80034 18920
rect 80074 18880 80116 18920
rect 80156 18880 80198 18920
rect 80238 18880 80280 18920
rect 80320 18880 80329 18920
rect 95063 18880 95072 18920
rect 95112 18880 95154 18920
rect 95194 18880 95236 18920
rect 95276 18880 95318 18920
rect 95358 18880 95400 18920
rect 95440 18880 95449 18920
rect 26467 18712 26476 18752
rect 26516 18712 32780 18752
rect 32740 18668 32780 18712
rect 21091 18628 21100 18668
rect 21140 18628 22444 18668
rect 22484 18628 23960 18668
rect 26083 18628 26092 18668
rect 26132 18628 27340 18668
rect 27380 18628 27389 18668
rect 32740 18628 36844 18668
rect 36884 18628 37228 18668
rect 37268 18628 37277 18668
rect 23920 18584 23960 18628
rect 23920 18544 26420 18584
rect 27427 18544 27436 18584
rect 27476 18544 28396 18584
rect 28436 18544 28445 18584
rect 26380 18500 26420 18544
rect 22723 18460 22732 18500
rect 22772 18460 26188 18500
rect 26228 18460 26237 18500
rect 26371 18460 26380 18500
rect 26420 18460 39052 18500
rect 39092 18460 39101 18500
rect 22435 18292 22444 18332
rect 22484 18292 22636 18332
rect 22676 18292 26476 18332
rect 26516 18292 26525 18332
rect 0 18248 80 18268
rect 0 18208 652 18248
rect 692 18208 701 18248
rect 0 18188 80 18208
rect 3103 18124 3112 18164
rect 3152 18124 3194 18164
rect 3234 18124 3276 18164
rect 3316 18124 3358 18164
rect 3398 18124 3440 18164
rect 3480 18124 3489 18164
rect 18223 18124 18232 18164
rect 18272 18124 18314 18164
rect 18354 18124 18396 18164
rect 18436 18124 18478 18164
rect 18518 18124 18560 18164
rect 18600 18124 18609 18164
rect 33343 18124 33352 18164
rect 33392 18124 33434 18164
rect 33474 18124 33516 18164
rect 33556 18124 33598 18164
rect 33638 18124 33680 18164
rect 33720 18124 33729 18164
rect 48463 18124 48472 18164
rect 48512 18124 48554 18164
rect 48594 18124 48636 18164
rect 48676 18124 48718 18164
rect 48758 18124 48800 18164
rect 48840 18124 48849 18164
rect 63583 18124 63592 18164
rect 63632 18124 63674 18164
rect 63714 18124 63756 18164
rect 63796 18124 63838 18164
rect 63878 18124 63920 18164
rect 63960 18124 63969 18164
rect 78703 18124 78712 18164
rect 78752 18124 78794 18164
rect 78834 18124 78876 18164
rect 78916 18124 78958 18164
rect 78998 18124 79040 18164
rect 79080 18124 79089 18164
rect 93823 18124 93832 18164
rect 93872 18124 93914 18164
rect 93954 18124 93996 18164
rect 94036 18124 94078 18164
rect 94118 18124 94160 18164
rect 94200 18124 94209 18164
rect 21379 17956 21388 17996
rect 21428 17956 22060 17996
rect 22100 17956 22252 17996
rect 22292 17956 22301 17996
rect 23920 17788 31372 17828
rect 31412 17788 31421 17828
rect 23920 17744 23960 17788
rect 16195 17704 16204 17744
rect 16244 17704 17644 17744
rect 17684 17704 17693 17744
rect 19363 17704 19372 17744
rect 19412 17704 22732 17744
rect 22772 17704 22781 17744
rect 22915 17704 22924 17744
rect 22964 17704 23960 17744
rect 26275 17704 26284 17744
rect 26324 17704 26764 17744
rect 26804 17704 26813 17744
rect 28003 17704 28012 17744
rect 28052 17704 32620 17744
rect 32660 17704 32669 17744
rect 33091 17704 33100 17744
rect 33140 17704 33676 17744
rect 33716 17704 33725 17744
rect 22243 17620 22252 17660
rect 22292 17620 22828 17660
rect 22868 17620 22877 17660
rect 28195 17620 28204 17660
rect 28244 17620 29164 17660
rect 29204 17620 29213 17660
rect 33763 17620 33772 17660
rect 33812 17620 34252 17660
rect 34292 17620 34301 17660
rect 0 17408 80 17428
rect 0 17368 652 17408
rect 692 17368 701 17408
rect 4343 17368 4352 17408
rect 4392 17368 4434 17408
rect 4474 17368 4516 17408
rect 4556 17368 4598 17408
rect 4638 17368 4680 17408
rect 4720 17368 4729 17408
rect 19463 17368 19472 17408
rect 19512 17368 19554 17408
rect 19594 17368 19636 17408
rect 19676 17368 19718 17408
rect 19758 17368 19800 17408
rect 19840 17368 19849 17408
rect 34583 17368 34592 17408
rect 34632 17368 34674 17408
rect 34714 17368 34756 17408
rect 34796 17368 34838 17408
rect 34878 17368 34920 17408
rect 34960 17368 34969 17408
rect 49703 17368 49712 17408
rect 49752 17368 49794 17408
rect 49834 17368 49876 17408
rect 49916 17368 49958 17408
rect 49998 17368 50040 17408
rect 50080 17368 50089 17408
rect 64823 17368 64832 17408
rect 64872 17368 64914 17408
rect 64954 17368 64996 17408
rect 65036 17368 65078 17408
rect 65118 17368 65160 17408
rect 65200 17368 65209 17408
rect 79943 17368 79952 17408
rect 79992 17368 80034 17408
rect 80074 17368 80116 17408
rect 80156 17368 80198 17408
rect 80238 17368 80280 17408
rect 80320 17368 80329 17408
rect 95063 17368 95072 17408
rect 95112 17368 95154 17408
rect 95194 17368 95236 17408
rect 95276 17368 95318 17408
rect 95358 17368 95400 17408
rect 95440 17368 95449 17408
rect 0 17348 80 17368
rect 31756 17116 37900 17156
rect 37940 17116 37949 17156
rect 31756 17072 31796 17116
rect 22243 17032 22252 17072
rect 22292 17032 22540 17072
rect 22580 17032 22589 17072
rect 27148 17032 31276 17072
rect 31316 17032 31756 17072
rect 31796 17032 31805 17072
rect 27148 16988 27188 17032
rect 23011 16948 23020 16988
rect 23060 16948 27148 16988
rect 27188 16948 27197 16988
rect 31171 16948 31180 16988
rect 31220 16948 34060 16988
rect 34100 16948 34109 16988
rect 3103 16612 3112 16652
rect 3152 16612 3194 16652
rect 3234 16612 3276 16652
rect 3316 16612 3358 16652
rect 3398 16612 3440 16652
rect 3480 16612 3489 16652
rect 18223 16612 18232 16652
rect 18272 16612 18314 16652
rect 18354 16612 18396 16652
rect 18436 16612 18478 16652
rect 18518 16612 18560 16652
rect 18600 16612 18609 16652
rect 33343 16612 33352 16652
rect 33392 16612 33434 16652
rect 33474 16612 33516 16652
rect 33556 16612 33598 16652
rect 33638 16612 33680 16652
rect 33720 16612 33729 16652
rect 48463 16612 48472 16652
rect 48512 16612 48554 16652
rect 48594 16612 48636 16652
rect 48676 16612 48718 16652
rect 48758 16612 48800 16652
rect 48840 16612 48849 16652
rect 63583 16612 63592 16652
rect 63632 16612 63674 16652
rect 63714 16612 63756 16652
rect 63796 16612 63838 16652
rect 63878 16612 63920 16652
rect 63960 16612 63969 16652
rect 78703 16612 78712 16652
rect 78752 16612 78794 16652
rect 78834 16612 78876 16652
rect 78916 16612 78958 16652
rect 78998 16612 79040 16652
rect 79080 16612 79089 16652
rect 93823 16612 93832 16652
rect 93872 16612 93914 16652
rect 93954 16612 93996 16652
rect 94036 16612 94078 16652
rect 94118 16612 94160 16652
rect 94200 16612 94209 16652
rect 0 16568 80 16588
rect 0 16528 652 16568
rect 692 16528 701 16568
rect 0 16508 80 16528
rect 30595 16360 30604 16400
rect 30644 16360 33196 16400
rect 33236 16360 33772 16400
rect 33812 16360 33821 16400
rect 34051 16276 34060 16316
rect 34100 16276 39244 16316
rect 39284 16276 40012 16316
rect 40052 16276 40061 16316
rect 37315 16192 37324 16232
rect 37364 16192 38572 16232
rect 38612 16192 38621 16232
rect 4343 15856 4352 15896
rect 4392 15856 4434 15896
rect 4474 15856 4516 15896
rect 4556 15856 4598 15896
rect 4638 15856 4680 15896
rect 4720 15856 4729 15896
rect 19463 15856 19472 15896
rect 19512 15856 19554 15896
rect 19594 15856 19636 15896
rect 19676 15856 19718 15896
rect 19758 15856 19800 15896
rect 19840 15856 19849 15896
rect 34583 15856 34592 15896
rect 34632 15856 34674 15896
rect 34714 15856 34756 15896
rect 34796 15856 34838 15896
rect 34878 15856 34920 15896
rect 34960 15856 34969 15896
rect 49703 15856 49712 15896
rect 49752 15856 49794 15896
rect 49834 15856 49876 15896
rect 49916 15856 49958 15896
rect 49998 15856 50040 15896
rect 50080 15856 50089 15896
rect 64823 15856 64832 15896
rect 64872 15856 64914 15896
rect 64954 15856 64996 15896
rect 65036 15856 65078 15896
rect 65118 15856 65160 15896
rect 65200 15856 65209 15896
rect 79943 15856 79952 15896
rect 79992 15856 80034 15896
rect 80074 15856 80116 15896
rect 80156 15856 80198 15896
rect 80238 15856 80280 15896
rect 80320 15856 80329 15896
rect 95063 15856 95072 15896
rect 95112 15856 95154 15896
rect 95194 15856 95236 15896
rect 95276 15856 95318 15896
rect 95358 15856 95400 15896
rect 95440 15856 95449 15896
rect 0 15728 80 15748
rect 0 15688 556 15728
rect 596 15688 605 15728
rect 17827 15688 17836 15728
rect 17876 15688 18220 15728
rect 18260 15688 18269 15728
rect 0 15668 80 15688
rect 16675 15520 16684 15560
rect 16724 15520 18988 15560
rect 19028 15520 20620 15560
rect 20660 15520 23788 15560
rect 23828 15520 23837 15560
rect 25027 15520 25036 15560
rect 25076 15520 27916 15560
rect 27956 15520 27965 15560
rect 28300 15520 33100 15560
rect 33140 15520 33149 15560
rect 28300 15476 28340 15520
rect 18403 15436 18412 15476
rect 18452 15436 28300 15476
rect 28340 15436 28349 15476
rect 18499 15352 18508 15392
rect 18548 15352 18892 15392
rect 18932 15352 18941 15392
rect 931 15268 940 15308
rect 980 15268 18700 15308
rect 18740 15268 18749 15308
rect 3103 15100 3112 15140
rect 3152 15100 3194 15140
rect 3234 15100 3276 15140
rect 3316 15100 3358 15140
rect 3398 15100 3440 15140
rect 3480 15100 3489 15140
rect 18223 15100 18232 15140
rect 18272 15100 18314 15140
rect 18354 15100 18396 15140
rect 18436 15100 18478 15140
rect 18518 15100 18560 15140
rect 18600 15100 18609 15140
rect 33343 15100 33352 15140
rect 33392 15100 33434 15140
rect 33474 15100 33516 15140
rect 33556 15100 33598 15140
rect 33638 15100 33680 15140
rect 33720 15100 33729 15140
rect 48463 15100 48472 15140
rect 48512 15100 48554 15140
rect 48594 15100 48636 15140
rect 48676 15100 48718 15140
rect 48758 15100 48800 15140
rect 48840 15100 48849 15140
rect 63583 15100 63592 15140
rect 63632 15100 63674 15140
rect 63714 15100 63756 15140
rect 63796 15100 63838 15140
rect 63878 15100 63920 15140
rect 63960 15100 63969 15140
rect 78703 15100 78712 15140
rect 78752 15100 78794 15140
rect 78834 15100 78876 15140
rect 78916 15100 78958 15140
rect 78998 15100 79040 15140
rect 79080 15100 79089 15140
rect 93823 15100 93832 15140
rect 93872 15100 93914 15140
rect 93954 15100 93996 15140
rect 94036 15100 94078 15140
rect 94118 15100 94160 15140
rect 94200 15100 94209 15140
rect 0 14888 80 14908
rect 0 14848 652 14888
rect 692 14848 701 14888
rect 0 14828 80 14848
rect 4343 14344 4352 14384
rect 4392 14344 4434 14384
rect 4474 14344 4516 14384
rect 4556 14344 4598 14384
rect 4638 14344 4680 14384
rect 4720 14344 4729 14384
rect 19463 14344 19472 14384
rect 19512 14344 19554 14384
rect 19594 14344 19636 14384
rect 19676 14344 19718 14384
rect 19758 14344 19800 14384
rect 19840 14344 19849 14384
rect 34583 14344 34592 14384
rect 34632 14344 34674 14384
rect 34714 14344 34756 14384
rect 34796 14344 34838 14384
rect 34878 14344 34920 14384
rect 34960 14344 34969 14384
rect 49703 14344 49712 14384
rect 49752 14344 49794 14384
rect 49834 14344 49876 14384
rect 49916 14344 49958 14384
rect 49998 14344 50040 14384
rect 50080 14344 50089 14384
rect 64823 14344 64832 14384
rect 64872 14344 64914 14384
rect 64954 14344 64996 14384
rect 65036 14344 65078 14384
rect 65118 14344 65160 14384
rect 65200 14344 65209 14384
rect 79943 14344 79952 14384
rect 79992 14344 80034 14384
rect 80074 14344 80116 14384
rect 80156 14344 80198 14384
rect 80238 14344 80280 14384
rect 80320 14344 80329 14384
rect 95063 14344 95072 14384
rect 95112 14344 95154 14384
rect 95194 14344 95236 14384
rect 95276 14344 95318 14384
rect 95358 14344 95400 14384
rect 95440 14344 95449 14384
rect 0 14048 80 14068
rect 0 14008 652 14048
rect 692 14008 701 14048
rect 0 13988 80 14008
rect 3103 13588 3112 13628
rect 3152 13588 3194 13628
rect 3234 13588 3276 13628
rect 3316 13588 3358 13628
rect 3398 13588 3440 13628
rect 3480 13588 3489 13628
rect 18223 13588 18232 13628
rect 18272 13588 18314 13628
rect 18354 13588 18396 13628
rect 18436 13588 18478 13628
rect 18518 13588 18560 13628
rect 18600 13588 18609 13628
rect 33343 13588 33352 13628
rect 33392 13588 33434 13628
rect 33474 13588 33516 13628
rect 33556 13588 33598 13628
rect 33638 13588 33680 13628
rect 33720 13588 33729 13628
rect 48463 13588 48472 13628
rect 48512 13588 48554 13628
rect 48594 13588 48636 13628
rect 48676 13588 48718 13628
rect 48758 13588 48800 13628
rect 48840 13588 48849 13628
rect 63583 13588 63592 13628
rect 63632 13588 63674 13628
rect 63714 13588 63756 13628
rect 63796 13588 63838 13628
rect 63878 13588 63920 13628
rect 63960 13588 63969 13628
rect 78703 13588 78712 13628
rect 78752 13588 78794 13628
rect 78834 13588 78876 13628
rect 78916 13588 78958 13628
rect 78998 13588 79040 13628
rect 79080 13588 79089 13628
rect 93823 13588 93832 13628
rect 93872 13588 93914 13628
rect 93954 13588 93996 13628
rect 94036 13588 94078 13628
rect 94118 13588 94160 13628
rect 94200 13588 94209 13628
rect 0 13208 80 13228
rect 0 13168 652 13208
rect 692 13168 701 13208
rect 26947 13168 26956 13208
rect 26996 13168 33196 13208
rect 33236 13168 34156 13208
rect 34196 13168 34205 13208
rect 0 13148 80 13168
rect 835 13000 844 13040
rect 884 13000 33004 13040
rect 33044 13000 33053 13040
rect 4343 12832 4352 12872
rect 4392 12832 4434 12872
rect 4474 12832 4516 12872
rect 4556 12832 4598 12872
rect 4638 12832 4680 12872
rect 4720 12832 4729 12872
rect 19463 12832 19472 12872
rect 19512 12832 19554 12872
rect 19594 12832 19636 12872
rect 19676 12832 19718 12872
rect 19758 12832 19800 12872
rect 19840 12832 19849 12872
rect 34583 12832 34592 12872
rect 34632 12832 34674 12872
rect 34714 12832 34756 12872
rect 34796 12832 34838 12872
rect 34878 12832 34920 12872
rect 34960 12832 34969 12872
rect 49703 12832 49712 12872
rect 49752 12832 49794 12872
rect 49834 12832 49876 12872
rect 49916 12832 49958 12872
rect 49998 12832 50040 12872
rect 50080 12832 50089 12872
rect 64823 12832 64832 12872
rect 64872 12832 64914 12872
rect 64954 12832 64996 12872
rect 65036 12832 65078 12872
rect 65118 12832 65160 12872
rect 65200 12832 65209 12872
rect 79943 12832 79952 12872
rect 79992 12832 80034 12872
rect 80074 12832 80116 12872
rect 80156 12832 80198 12872
rect 80238 12832 80280 12872
rect 80320 12832 80329 12872
rect 95063 12832 95072 12872
rect 95112 12832 95154 12872
rect 95194 12832 95236 12872
rect 95276 12832 95318 12872
rect 95358 12832 95400 12872
rect 95440 12832 95449 12872
rect 26851 12748 26860 12788
rect 26900 12748 27820 12788
rect 27860 12748 27869 12788
rect 26563 12664 26572 12704
rect 26612 12664 26956 12704
rect 26996 12664 27005 12704
rect 26467 12580 26476 12620
rect 26516 12580 27244 12620
rect 27284 12580 27293 12620
rect 15811 12496 15820 12536
rect 15860 12496 18124 12536
rect 18164 12496 23020 12536
rect 23060 12496 23069 12536
rect 27427 12412 27436 12452
rect 27476 12412 28012 12452
rect 28052 12412 28061 12452
rect 0 12368 80 12388
rect 0 12328 652 12368
rect 692 12328 701 12368
rect 0 12308 80 12328
rect 20131 12244 20140 12284
rect 20180 12244 26764 12284
rect 26804 12244 26813 12284
rect 27235 12244 27244 12284
rect 27284 12244 27293 12284
rect 27244 12200 27284 12244
rect 739 12160 748 12200
rect 788 12160 27284 12200
rect 3103 12076 3112 12116
rect 3152 12076 3194 12116
rect 3234 12076 3276 12116
rect 3316 12076 3358 12116
rect 3398 12076 3440 12116
rect 3480 12076 3489 12116
rect 18223 12076 18232 12116
rect 18272 12076 18314 12116
rect 18354 12076 18396 12116
rect 18436 12076 18478 12116
rect 18518 12076 18560 12116
rect 18600 12076 18609 12116
rect 33343 12076 33352 12116
rect 33392 12076 33434 12116
rect 33474 12076 33516 12116
rect 33556 12076 33598 12116
rect 33638 12076 33680 12116
rect 33720 12076 33729 12116
rect 48463 12076 48472 12116
rect 48512 12076 48554 12116
rect 48594 12076 48636 12116
rect 48676 12076 48718 12116
rect 48758 12076 48800 12116
rect 48840 12076 48849 12116
rect 63583 12076 63592 12116
rect 63632 12076 63674 12116
rect 63714 12076 63756 12116
rect 63796 12076 63838 12116
rect 63878 12076 63920 12116
rect 63960 12076 63969 12116
rect 78703 12076 78712 12116
rect 78752 12076 78794 12116
rect 78834 12076 78876 12116
rect 78916 12076 78958 12116
rect 78998 12076 79040 12116
rect 79080 12076 79089 12116
rect 93823 12076 93832 12116
rect 93872 12076 93914 12116
rect 93954 12076 93996 12116
rect 94036 12076 94078 12116
rect 94118 12076 94160 12116
rect 94200 12076 94209 12116
rect 1027 11992 1036 12032
rect 1076 11992 27820 12032
rect 27860 11992 27869 12032
rect 24931 11908 24940 11948
rect 24980 11908 26380 11948
rect 26420 11908 26429 11948
rect 0 11528 80 11548
rect 0 11488 652 11528
rect 692 11488 701 11528
rect 0 11468 80 11488
rect 4343 11320 4352 11360
rect 4392 11320 4434 11360
rect 4474 11320 4516 11360
rect 4556 11320 4598 11360
rect 4638 11320 4680 11360
rect 4720 11320 4729 11360
rect 19463 11320 19472 11360
rect 19512 11320 19554 11360
rect 19594 11320 19636 11360
rect 19676 11320 19718 11360
rect 19758 11320 19800 11360
rect 19840 11320 19849 11360
rect 34583 11320 34592 11360
rect 34632 11320 34674 11360
rect 34714 11320 34756 11360
rect 34796 11320 34838 11360
rect 34878 11320 34920 11360
rect 34960 11320 34969 11360
rect 49703 11320 49712 11360
rect 49752 11320 49794 11360
rect 49834 11320 49876 11360
rect 49916 11320 49958 11360
rect 49998 11320 50040 11360
rect 50080 11320 50089 11360
rect 64823 11320 64832 11360
rect 64872 11320 64914 11360
rect 64954 11320 64996 11360
rect 65036 11320 65078 11360
rect 65118 11320 65160 11360
rect 65200 11320 65209 11360
rect 79943 11320 79952 11360
rect 79992 11320 80034 11360
rect 80074 11320 80116 11360
rect 80156 11320 80198 11360
rect 80238 11320 80280 11360
rect 80320 11320 80329 11360
rect 95063 11320 95072 11360
rect 95112 11320 95154 11360
rect 95194 11320 95236 11360
rect 95276 11320 95318 11360
rect 95358 11320 95400 11360
rect 95440 11320 95449 11360
rect 835 10900 844 10940
rect 884 10900 18028 10940
rect 18068 10900 18077 10940
rect 643 10732 652 10772
rect 692 10732 701 10772
rect 0 10688 80 10708
rect 652 10688 692 10732
rect 0 10648 692 10688
rect 0 10628 80 10648
rect 3103 10564 3112 10604
rect 3152 10564 3194 10604
rect 3234 10564 3276 10604
rect 3316 10564 3358 10604
rect 3398 10564 3440 10604
rect 3480 10564 3489 10604
rect 18223 10564 18232 10604
rect 18272 10564 18314 10604
rect 18354 10564 18396 10604
rect 18436 10564 18478 10604
rect 18518 10564 18560 10604
rect 18600 10564 18609 10604
rect 33343 10564 33352 10604
rect 33392 10564 33434 10604
rect 33474 10564 33516 10604
rect 33556 10564 33598 10604
rect 33638 10564 33680 10604
rect 33720 10564 33729 10604
rect 48463 10564 48472 10604
rect 48512 10564 48554 10604
rect 48594 10564 48636 10604
rect 48676 10564 48718 10604
rect 48758 10564 48800 10604
rect 48840 10564 48849 10604
rect 63583 10564 63592 10604
rect 63632 10564 63674 10604
rect 63714 10564 63756 10604
rect 63796 10564 63838 10604
rect 63878 10564 63920 10604
rect 63960 10564 63969 10604
rect 78703 10564 78712 10604
rect 78752 10564 78794 10604
rect 78834 10564 78876 10604
rect 78916 10564 78958 10604
rect 78998 10564 79040 10604
rect 79080 10564 79089 10604
rect 93823 10564 93832 10604
rect 93872 10564 93914 10604
rect 93954 10564 93996 10604
rect 94036 10564 94078 10604
rect 94118 10564 94160 10604
rect 94200 10564 94209 10604
rect 835 10228 844 10268
rect 884 10228 36748 10268
rect 36788 10228 36797 10268
rect 0 9848 80 9868
rect 0 9808 652 9848
rect 692 9808 701 9848
rect 4343 9808 4352 9848
rect 4392 9808 4434 9848
rect 4474 9808 4516 9848
rect 4556 9808 4598 9848
rect 4638 9808 4680 9848
rect 4720 9808 4729 9848
rect 19463 9808 19472 9848
rect 19512 9808 19554 9848
rect 19594 9808 19636 9848
rect 19676 9808 19718 9848
rect 19758 9808 19800 9848
rect 19840 9808 19849 9848
rect 34583 9808 34592 9848
rect 34632 9808 34674 9848
rect 34714 9808 34756 9848
rect 34796 9808 34838 9848
rect 34878 9808 34920 9848
rect 34960 9808 34969 9848
rect 49703 9808 49712 9848
rect 49752 9808 49794 9848
rect 49834 9808 49876 9848
rect 49916 9808 49958 9848
rect 49998 9808 50040 9848
rect 50080 9808 50089 9848
rect 64823 9808 64832 9848
rect 64872 9808 64914 9848
rect 64954 9808 64996 9848
rect 65036 9808 65078 9848
rect 65118 9808 65160 9848
rect 65200 9808 65209 9848
rect 79943 9808 79952 9848
rect 79992 9808 80034 9848
rect 80074 9808 80116 9848
rect 80156 9808 80198 9848
rect 80238 9808 80280 9848
rect 80320 9808 80329 9848
rect 95063 9808 95072 9848
rect 95112 9808 95154 9848
rect 95194 9808 95236 9848
rect 95276 9808 95318 9848
rect 95358 9808 95400 9848
rect 95440 9808 95449 9848
rect 0 9788 80 9808
rect 835 9388 844 9428
rect 884 9388 27052 9428
rect 27092 9388 27101 9428
rect 3103 9052 3112 9092
rect 3152 9052 3194 9092
rect 3234 9052 3276 9092
rect 3316 9052 3358 9092
rect 3398 9052 3440 9092
rect 3480 9052 3489 9092
rect 18223 9052 18232 9092
rect 18272 9052 18314 9092
rect 18354 9052 18396 9092
rect 18436 9052 18478 9092
rect 18518 9052 18560 9092
rect 18600 9052 18609 9092
rect 33343 9052 33352 9092
rect 33392 9052 33434 9092
rect 33474 9052 33516 9092
rect 33556 9052 33598 9092
rect 33638 9052 33680 9092
rect 33720 9052 33729 9092
rect 48463 9052 48472 9092
rect 48512 9052 48554 9092
rect 48594 9052 48636 9092
rect 48676 9052 48718 9092
rect 48758 9052 48800 9092
rect 48840 9052 48849 9092
rect 63583 9052 63592 9092
rect 63632 9052 63674 9092
rect 63714 9052 63756 9092
rect 63796 9052 63838 9092
rect 63878 9052 63920 9092
rect 63960 9052 63969 9092
rect 78703 9052 78712 9092
rect 78752 9052 78794 9092
rect 78834 9052 78876 9092
rect 78916 9052 78958 9092
rect 78998 9052 79040 9092
rect 79080 9052 79089 9092
rect 93823 9052 93832 9092
rect 93872 9052 93914 9092
rect 93954 9052 93996 9092
rect 94036 9052 94078 9092
rect 94118 9052 94160 9092
rect 94200 9052 94209 9092
rect 0 9008 80 9028
rect 0 8968 652 9008
rect 692 8968 701 9008
rect 0 8948 80 8968
rect 4343 8296 4352 8336
rect 4392 8296 4434 8336
rect 4474 8296 4516 8336
rect 4556 8296 4598 8336
rect 4638 8296 4680 8336
rect 4720 8296 4729 8336
rect 19463 8296 19472 8336
rect 19512 8296 19554 8336
rect 19594 8296 19636 8336
rect 19676 8296 19718 8336
rect 19758 8296 19800 8336
rect 19840 8296 19849 8336
rect 34583 8296 34592 8336
rect 34632 8296 34674 8336
rect 34714 8296 34756 8336
rect 34796 8296 34838 8336
rect 34878 8296 34920 8336
rect 34960 8296 34969 8336
rect 49703 8296 49712 8336
rect 49752 8296 49794 8336
rect 49834 8296 49876 8336
rect 49916 8296 49958 8336
rect 49998 8296 50040 8336
rect 50080 8296 50089 8336
rect 64823 8296 64832 8336
rect 64872 8296 64914 8336
rect 64954 8296 64996 8336
rect 65036 8296 65078 8336
rect 65118 8296 65160 8336
rect 65200 8296 65209 8336
rect 79943 8296 79952 8336
rect 79992 8296 80034 8336
rect 80074 8296 80116 8336
rect 80156 8296 80198 8336
rect 80238 8296 80280 8336
rect 80320 8296 80329 8336
rect 95063 8296 95072 8336
rect 95112 8296 95154 8336
rect 95194 8296 95236 8336
rect 95276 8296 95318 8336
rect 95358 8296 95400 8336
rect 95440 8296 95449 8336
rect 0 8168 80 8188
rect 0 8128 652 8168
rect 692 8128 701 8168
rect 0 8108 80 8128
rect 3103 7540 3112 7580
rect 3152 7540 3194 7580
rect 3234 7540 3276 7580
rect 3316 7540 3358 7580
rect 3398 7540 3440 7580
rect 3480 7540 3489 7580
rect 18223 7540 18232 7580
rect 18272 7540 18314 7580
rect 18354 7540 18396 7580
rect 18436 7540 18478 7580
rect 18518 7540 18560 7580
rect 18600 7540 18609 7580
rect 33343 7540 33352 7580
rect 33392 7540 33434 7580
rect 33474 7540 33516 7580
rect 33556 7540 33598 7580
rect 33638 7540 33680 7580
rect 33720 7540 33729 7580
rect 48463 7540 48472 7580
rect 48512 7540 48554 7580
rect 48594 7540 48636 7580
rect 48676 7540 48718 7580
rect 48758 7540 48800 7580
rect 48840 7540 48849 7580
rect 63583 7540 63592 7580
rect 63632 7540 63674 7580
rect 63714 7540 63756 7580
rect 63796 7540 63838 7580
rect 63878 7540 63920 7580
rect 63960 7540 63969 7580
rect 78703 7540 78712 7580
rect 78752 7540 78794 7580
rect 78834 7540 78876 7580
rect 78916 7540 78958 7580
rect 78998 7540 79040 7580
rect 79080 7540 79089 7580
rect 93823 7540 93832 7580
rect 93872 7540 93914 7580
rect 93954 7540 93996 7580
rect 94036 7540 94078 7580
rect 94118 7540 94160 7580
rect 94200 7540 94209 7580
rect 0 7328 80 7348
rect 0 7288 652 7328
rect 692 7288 701 7328
rect 0 7268 80 7288
rect 835 7204 844 7244
rect 884 7204 34252 7244
rect 34292 7204 34301 7244
rect 4343 6784 4352 6824
rect 4392 6784 4434 6824
rect 4474 6784 4516 6824
rect 4556 6784 4598 6824
rect 4638 6784 4680 6824
rect 4720 6784 4729 6824
rect 19463 6784 19472 6824
rect 19512 6784 19554 6824
rect 19594 6784 19636 6824
rect 19676 6784 19718 6824
rect 19758 6784 19800 6824
rect 19840 6784 19849 6824
rect 34583 6784 34592 6824
rect 34632 6784 34674 6824
rect 34714 6784 34756 6824
rect 34796 6784 34838 6824
rect 34878 6784 34920 6824
rect 34960 6784 34969 6824
rect 49703 6784 49712 6824
rect 49752 6784 49794 6824
rect 49834 6784 49876 6824
rect 49916 6784 49958 6824
rect 49998 6784 50040 6824
rect 50080 6784 50089 6824
rect 64823 6784 64832 6824
rect 64872 6784 64914 6824
rect 64954 6784 64996 6824
rect 65036 6784 65078 6824
rect 65118 6784 65160 6824
rect 65200 6784 65209 6824
rect 79943 6784 79952 6824
rect 79992 6784 80034 6824
rect 80074 6784 80116 6824
rect 80156 6784 80198 6824
rect 80238 6784 80280 6824
rect 80320 6784 80329 6824
rect 95063 6784 95072 6824
rect 95112 6784 95154 6824
rect 95194 6784 95236 6824
rect 95276 6784 95318 6824
rect 95358 6784 95400 6824
rect 95440 6784 95449 6824
rect 0 6488 80 6508
rect 0 6448 652 6488
rect 692 6448 701 6488
rect 0 6428 80 6448
rect 3103 6028 3112 6068
rect 3152 6028 3194 6068
rect 3234 6028 3276 6068
rect 3316 6028 3358 6068
rect 3398 6028 3440 6068
rect 3480 6028 3489 6068
rect 18223 6028 18232 6068
rect 18272 6028 18314 6068
rect 18354 6028 18396 6068
rect 18436 6028 18478 6068
rect 18518 6028 18560 6068
rect 18600 6028 18609 6068
rect 33343 6028 33352 6068
rect 33392 6028 33434 6068
rect 33474 6028 33516 6068
rect 33556 6028 33598 6068
rect 33638 6028 33680 6068
rect 33720 6028 33729 6068
rect 48463 6028 48472 6068
rect 48512 6028 48554 6068
rect 48594 6028 48636 6068
rect 48676 6028 48718 6068
rect 48758 6028 48800 6068
rect 48840 6028 48849 6068
rect 63583 6028 63592 6068
rect 63632 6028 63674 6068
rect 63714 6028 63756 6068
rect 63796 6028 63838 6068
rect 63878 6028 63920 6068
rect 63960 6028 63969 6068
rect 78703 6028 78712 6068
rect 78752 6028 78794 6068
rect 78834 6028 78876 6068
rect 78916 6028 78958 6068
rect 78998 6028 79040 6068
rect 79080 6028 79089 6068
rect 93823 6028 93832 6068
rect 93872 6028 93914 6068
rect 93954 6028 93996 6068
rect 94036 6028 94078 6068
rect 94118 6028 94160 6068
rect 94200 6028 94209 6068
rect 835 5692 844 5732
rect 884 5692 18700 5732
rect 18740 5692 18749 5732
rect 0 5648 80 5668
rect 0 5608 652 5648
rect 692 5608 701 5648
rect 0 5588 80 5608
rect 4343 5272 4352 5312
rect 4392 5272 4434 5312
rect 4474 5272 4516 5312
rect 4556 5272 4598 5312
rect 4638 5272 4680 5312
rect 4720 5272 4729 5312
rect 19463 5272 19472 5312
rect 19512 5272 19554 5312
rect 19594 5272 19636 5312
rect 19676 5272 19718 5312
rect 19758 5272 19800 5312
rect 19840 5272 19849 5312
rect 34583 5272 34592 5312
rect 34632 5272 34674 5312
rect 34714 5272 34756 5312
rect 34796 5272 34838 5312
rect 34878 5272 34920 5312
rect 34960 5272 34969 5312
rect 49703 5272 49712 5312
rect 49752 5272 49794 5312
rect 49834 5272 49876 5312
rect 49916 5272 49958 5312
rect 49998 5272 50040 5312
rect 50080 5272 50089 5312
rect 64823 5272 64832 5312
rect 64872 5272 64914 5312
rect 64954 5272 64996 5312
rect 65036 5272 65078 5312
rect 65118 5272 65160 5312
rect 65200 5272 65209 5312
rect 79943 5272 79952 5312
rect 79992 5272 80034 5312
rect 80074 5272 80116 5312
rect 80156 5272 80198 5312
rect 80238 5272 80280 5312
rect 80320 5272 80329 5312
rect 95063 5272 95072 5312
rect 95112 5272 95154 5312
rect 95194 5272 95236 5312
rect 95276 5272 95318 5312
rect 95358 5272 95400 5312
rect 95440 5272 95449 5312
rect 835 4852 844 4892
rect 884 4852 34348 4892
rect 34388 4852 34397 4892
rect 0 4808 80 4828
rect 0 4768 652 4808
rect 692 4768 701 4808
rect 0 4748 80 4768
rect 3103 4516 3112 4556
rect 3152 4516 3194 4556
rect 3234 4516 3276 4556
rect 3316 4516 3358 4556
rect 3398 4516 3440 4556
rect 3480 4516 3489 4556
rect 18223 4516 18232 4556
rect 18272 4516 18314 4556
rect 18354 4516 18396 4556
rect 18436 4516 18478 4556
rect 18518 4516 18560 4556
rect 18600 4516 18609 4556
rect 33343 4516 33352 4556
rect 33392 4516 33434 4556
rect 33474 4516 33516 4556
rect 33556 4516 33598 4556
rect 33638 4516 33680 4556
rect 33720 4516 33729 4556
rect 48463 4516 48472 4556
rect 48512 4516 48554 4556
rect 48594 4516 48636 4556
rect 48676 4516 48718 4556
rect 48758 4516 48800 4556
rect 48840 4516 48849 4556
rect 63583 4516 63592 4556
rect 63632 4516 63674 4556
rect 63714 4516 63756 4556
rect 63796 4516 63838 4556
rect 63878 4516 63920 4556
rect 63960 4516 63969 4556
rect 78703 4516 78712 4556
rect 78752 4516 78794 4556
rect 78834 4516 78876 4556
rect 78916 4516 78958 4556
rect 78998 4516 79040 4556
rect 79080 4516 79089 4556
rect 93823 4516 93832 4556
rect 93872 4516 93914 4556
rect 93954 4516 93996 4556
rect 94036 4516 94078 4556
rect 94118 4516 94160 4556
rect 94200 4516 94209 4556
rect 835 4180 844 4220
rect 884 4180 34444 4220
rect 34484 4180 34493 4220
rect 0 3968 80 3988
rect 0 3928 652 3968
rect 692 3928 701 3968
rect 0 3908 80 3928
rect 4343 3760 4352 3800
rect 4392 3760 4434 3800
rect 4474 3760 4516 3800
rect 4556 3760 4598 3800
rect 4638 3760 4680 3800
rect 4720 3760 4729 3800
rect 19463 3760 19472 3800
rect 19512 3760 19554 3800
rect 19594 3760 19636 3800
rect 19676 3760 19718 3800
rect 19758 3760 19800 3800
rect 19840 3760 19849 3800
rect 34583 3760 34592 3800
rect 34632 3760 34674 3800
rect 34714 3760 34756 3800
rect 34796 3760 34838 3800
rect 34878 3760 34920 3800
rect 34960 3760 34969 3800
rect 49703 3760 49712 3800
rect 49752 3760 49794 3800
rect 49834 3760 49876 3800
rect 49916 3760 49958 3800
rect 49998 3760 50040 3800
rect 50080 3760 50089 3800
rect 64823 3760 64832 3800
rect 64872 3760 64914 3800
rect 64954 3760 64996 3800
rect 65036 3760 65078 3800
rect 65118 3760 65160 3800
rect 65200 3760 65209 3800
rect 79943 3760 79952 3800
rect 79992 3760 80034 3800
rect 80074 3760 80116 3800
rect 80156 3760 80198 3800
rect 80238 3760 80280 3800
rect 80320 3760 80329 3800
rect 95063 3760 95072 3800
rect 95112 3760 95154 3800
rect 95194 3760 95236 3800
rect 95276 3760 95318 3800
rect 95358 3760 95400 3800
rect 95440 3760 95449 3800
rect 643 3172 652 3212
rect 692 3172 701 3212
rect 0 3128 80 3148
rect 652 3128 692 3172
rect 0 3088 692 3128
rect 0 3068 80 3088
rect 3103 3004 3112 3044
rect 3152 3004 3194 3044
rect 3234 3004 3276 3044
rect 3316 3004 3358 3044
rect 3398 3004 3440 3044
rect 3480 3004 3489 3044
rect 18223 3004 18232 3044
rect 18272 3004 18314 3044
rect 18354 3004 18396 3044
rect 18436 3004 18478 3044
rect 18518 3004 18560 3044
rect 18600 3004 18609 3044
rect 33343 3004 33352 3044
rect 33392 3004 33434 3044
rect 33474 3004 33516 3044
rect 33556 3004 33598 3044
rect 33638 3004 33680 3044
rect 33720 3004 33729 3044
rect 48463 3004 48472 3044
rect 48512 3004 48554 3044
rect 48594 3004 48636 3044
rect 48676 3004 48718 3044
rect 48758 3004 48800 3044
rect 48840 3004 48849 3044
rect 63583 3004 63592 3044
rect 63632 3004 63674 3044
rect 63714 3004 63756 3044
rect 63796 3004 63838 3044
rect 63878 3004 63920 3044
rect 63960 3004 63969 3044
rect 78703 3004 78712 3044
rect 78752 3004 78794 3044
rect 78834 3004 78876 3044
rect 78916 3004 78958 3044
rect 78998 3004 79040 3044
rect 79080 3004 79089 3044
rect 93823 3004 93832 3044
rect 93872 3004 93914 3044
rect 93954 3004 93996 3044
rect 94036 3004 94078 3044
rect 94118 3004 94160 3044
rect 94200 3004 94209 3044
rect 0 2288 80 2308
rect 0 2248 652 2288
rect 692 2248 701 2288
rect 4343 2248 4352 2288
rect 4392 2248 4434 2288
rect 4474 2248 4516 2288
rect 4556 2248 4598 2288
rect 4638 2248 4680 2288
rect 4720 2248 4729 2288
rect 19463 2248 19472 2288
rect 19512 2248 19554 2288
rect 19594 2248 19636 2288
rect 19676 2248 19718 2288
rect 19758 2248 19800 2288
rect 19840 2248 19849 2288
rect 34583 2248 34592 2288
rect 34632 2248 34674 2288
rect 34714 2248 34756 2288
rect 34796 2248 34838 2288
rect 34878 2248 34920 2288
rect 34960 2248 34969 2288
rect 49703 2248 49712 2288
rect 49752 2248 49794 2288
rect 49834 2248 49876 2288
rect 49916 2248 49958 2288
rect 49998 2248 50040 2288
rect 50080 2248 50089 2288
rect 64823 2248 64832 2288
rect 64872 2248 64914 2288
rect 64954 2248 64996 2288
rect 65036 2248 65078 2288
rect 65118 2248 65160 2288
rect 65200 2248 65209 2288
rect 79943 2248 79952 2288
rect 79992 2248 80034 2288
rect 80074 2248 80116 2288
rect 80156 2248 80198 2288
rect 80238 2248 80280 2288
rect 80320 2248 80329 2288
rect 95063 2248 95072 2288
rect 95112 2248 95154 2288
rect 95194 2248 95236 2288
rect 95276 2248 95318 2288
rect 95358 2248 95400 2288
rect 95440 2248 95449 2288
rect 0 2228 80 2248
rect 3103 1492 3112 1532
rect 3152 1492 3194 1532
rect 3234 1492 3276 1532
rect 3316 1492 3358 1532
rect 3398 1492 3440 1532
rect 3480 1492 3489 1532
rect 18223 1492 18232 1532
rect 18272 1492 18314 1532
rect 18354 1492 18396 1532
rect 18436 1492 18478 1532
rect 18518 1492 18560 1532
rect 18600 1492 18609 1532
rect 33343 1492 33352 1532
rect 33392 1492 33434 1532
rect 33474 1492 33516 1532
rect 33556 1492 33598 1532
rect 33638 1492 33680 1532
rect 33720 1492 33729 1532
rect 48463 1492 48472 1532
rect 48512 1492 48554 1532
rect 48594 1492 48636 1532
rect 48676 1492 48718 1532
rect 48758 1492 48800 1532
rect 48840 1492 48849 1532
rect 63583 1492 63592 1532
rect 63632 1492 63674 1532
rect 63714 1492 63756 1532
rect 63796 1492 63838 1532
rect 63878 1492 63920 1532
rect 63960 1492 63969 1532
rect 78703 1492 78712 1532
rect 78752 1492 78794 1532
rect 78834 1492 78876 1532
rect 78916 1492 78958 1532
rect 78998 1492 79040 1532
rect 79080 1492 79089 1532
rect 93823 1492 93832 1532
rect 93872 1492 93914 1532
rect 93954 1492 93996 1532
rect 94036 1492 94078 1532
rect 94118 1492 94160 1532
rect 94200 1492 94209 1532
rect 4343 736 4352 776
rect 4392 736 4434 776
rect 4474 736 4516 776
rect 4556 736 4598 776
rect 4638 736 4680 776
rect 4720 736 4729 776
rect 19463 736 19472 776
rect 19512 736 19554 776
rect 19594 736 19636 776
rect 19676 736 19718 776
rect 19758 736 19800 776
rect 19840 736 19849 776
rect 34583 736 34592 776
rect 34632 736 34674 776
rect 34714 736 34756 776
rect 34796 736 34838 776
rect 34878 736 34920 776
rect 34960 736 34969 776
rect 49703 736 49712 776
rect 49752 736 49794 776
rect 49834 736 49876 776
rect 49916 736 49958 776
rect 49998 736 50040 776
rect 50080 736 50089 776
rect 64823 736 64832 776
rect 64872 736 64914 776
rect 64954 736 64996 776
rect 65036 736 65078 776
rect 65118 736 65160 776
rect 65200 736 65209 776
rect 79943 736 79952 776
rect 79992 736 80034 776
rect 80074 736 80116 776
rect 80156 736 80198 776
rect 80238 736 80280 776
rect 80320 736 80329 776
rect 95063 736 95072 776
rect 95112 736 95154 776
rect 95194 736 95236 776
rect 95276 736 95318 776
rect 95358 736 95400 776
rect 95440 736 95449 776
<< via3 >>
rect 4352 38536 4392 38576
rect 4434 38536 4474 38576
rect 4516 38536 4556 38576
rect 4598 38536 4638 38576
rect 4680 38536 4720 38576
rect 19472 38536 19512 38576
rect 19554 38536 19594 38576
rect 19636 38536 19676 38576
rect 19718 38536 19758 38576
rect 19800 38536 19840 38576
rect 34592 38536 34632 38576
rect 34674 38536 34714 38576
rect 34756 38536 34796 38576
rect 34838 38536 34878 38576
rect 34920 38536 34960 38576
rect 49712 38536 49752 38576
rect 49794 38536 49834 38576
rect 49876 38536 49916 38576
rect 49958 38536 49998 38576
rect 50040 38536 50080 38576
rect 64832 38536 64872 38576
rect 64914 38536 64954 38576
rect 64996 38536 65036 38576
rect 65078 38536 65118 38576
rect 65160 38536 65200 38576
rect 79952 38536 79992 38576
rect 80034 38536 80074 38576
rect 80116 38536 80156 38576
rect 80198 38536 80238 38576
rect 80280 38536 80320 38576
rect 95072 38536 95112 38576
rect 95154 38536 95194 38576
rect 95236 38536 95276 38576
rect 95318 38536 95358 38576
rect 95400 38536 95440 38576
rect 3112 37780 3152 37820
rect 3194 37780 3234 37820
rect 3276 37780 3316 37820
rect 3358 37780 3398 37820
rect 3440 37780 3480 37820
rect 18232 37780 18272 37820
rect 18314 37780 18354 37820
rect 18396 37780 18436 37820
rect 18478 37780 18518 37820
rect 18560 37780 18600 37820
rect 33352 37780 33392 37820
rect 33434 37780 33474 37820
rect 33516 37780 33556 37820
rect 33598 37780 33638 37820
rect 33680 37780 33720 37820
rect 48472 37780 48512 37820
rect 48554 37780 48594 37820
rect 48636 37780 48676 37820
rect 48718 37780 48758 37820
rect 48800 37780 48840 37820
rect 63592 37780 63632 37820
rect 63674 37780 63714 37820
rect 63756 37780 63796 37820
rect 63838 37780 63878 37820
rect 63920 37780 63960 37820
rect 78712 37780 78752 37820
rect 78794 37780 78834 37820
rect 78876 37780 78916 37820
rect 78958 37780 78998 37820
rect 79040 37780 79080 37820
rect 93832 37780 93872 37820
rect 93914 37780 93954 37820
rect 93996 37780 94036 37820
rect 94078 37780 94118 37820
rect 94160 37780 94200 37820
rect 4352 37024 4392 37064
rect 4434 37024 4474 37064
rect 4516 37024 4556 37064
rect 4598 37024 4638 37064
rect 4680 37024 4720 37064
rect 19472 37024 19512 37064
rect 19554 37024 19594 37064
rect 19636 37024 19676 37064
rect 19718 37024 19758 37064
rect 19800 37024 19840 37064
rect 34592 37024 34632 37064
rect 34674 37024 34714 37064
rect 34756 37024 34796 37064
rect 34838 37024 34878 37064
rect 34920 37024 34960 37064
rect 49712 37024 49752 37064
rect 49794 37024 49834 37064
rect 49876 37024 49916 37064
rect 49958 37024 49998 37064
rect 50040 37024 50080 37064
rect 64832 37024 64872 37064
rect 64914 37024 64954 37064
rect 64996 37024 65036 37064
rect 65078 37024 65118 37064
rect 65160 37024 65200 37064
rect 79952 37024 79992 37064
rect 80034 37024 80074 37064
rect 80116 37024 80156 37064
rect 80198 37024 80238 37064
rect 80280 37024 80320 37064
rect 95072 37024 95112 37064
rect 95154 37024 95194 37064
rect 95236 37024 95276 37064
rect 95318 37024 95358 37064
rect 95400 37024 95440 37064
rect 3112 36268 3152 36308
rect 3194 36268 3234 36308
rect 3276 36268 3316 36308
rect 3358 36268 3398 36308
rect 3440 36268 3480 36308
rect 18232 36268 18272 36308
rect 18314 36268 18354 36308
rect 18396 36268 18436 36308
rect 18478 36268 18518 36308
rect 18560 36268 18600 36308
rect 33352 36268 33392 36308
rect 33434 36268 33474 36308
rect 33516 36268 33556 36308
rect 33598 36268 33638 36308
rect 33680 36268 33720 36308
rect 48472 36268 48512 36308
rect 48554 36268 48594 36308
rect 48636 36268 48676 36308
rect 48718 36268 48758 36308
rect 48800 36268 48840 36308
rect 63592 36268 63632 36308
rect 63674 36268 63714 36308
rect 63756 36268 63796 36308
rect 63838 36268 63878 36308
rect 63920 36268 63960 36308
rect 78712 36268 78752 36308
rect 78794 36268 78834 36308
rect 78876 36268 78916 36308
rect 78958 36268 78998 36308
rect 79040 36268 79080 36308
rect 93832 36268 93872 36308
rect 93914 36268 93954 36308
rect 93996 36268 94036 36308
rect 94078 36268 94118 36308
rect 94160 36268 94200 36308
rect 4352 35512 4392 35552
rect 4434 35512 4474 35552
rect 4516 35512 4556 35552
rect 4598 35512 4638 35552
rect 4680 35512 4720 35552
rect 19472 35512 19512 35552
rect 19554 35512 19594 35552
rect 19636 35512 19676 35552
rect 19718 35512 19758 35552
rect 19800 35512 19840 35552
rect 34592 35512 34632 35552
rect 34674 35512 34714 35552
rect 34756 35512 34796 35552
rect 34838 35512 34878 35552
rect 34920 35512 34960 35552
rect 49712 35512 49752 35552
rect 49794 35512 49834 35552
rect 49876 35512 49916 35552
rect 49958 35512 49998 35552
rect 50040 35512 50080 35552
rect 64832 35512 64872 35552
rect 64914 35512 64954 35552
rect 64996 35512 65036 35552
rect 65078 35512 65118 35552
rect 65160 35512 65200 35552
rect 79952 35512 79992 35552
rect 80034 35512 80074 35552
rect 80116 35512 80156 35552
rect 80198 35512 80238 35552
rect 80280 35512 80320 35552
rect 95072 35512 95112 35552
rect 95154 35512 95194 35552
rect 95236 35512 95276 35552
rect 95318 35512 95358 35552
rect 95400 35512 95440 35552
rect 3112 34756 3152 34796
rect 3194 34756 3234 34796
rect 3276 34756 3316 34796
rect 3358 34756 3398 34796
rect 3440 34756 3480 34796
rect 18232 34756 18272 34796
rect 18314 34756 18354 34796
rect 18396 34756 18436 34796
rect 18478 34756 18518 34796
rect 18560 34756 18600 34796
rect 33352 34756 33392 34796
rect 33434 34756 33474 34796
rect 33516 34756 33556 34796
rect 33598 34756 33638 34796
rect 33680 34756 33720 34796
rect 48472 34756 48512 34796
rect 48554 34756 48594 34796
rect 48636 34756 48676 34796
rect 48718 34756 48758 34796
rect 48800 34756 48840 34796
rect 63592 34756 63632 34796
rect 63674 34756 63714 34796
rect 63756 34756 63796 34796
rect 63838 34756 63878 34796
rect 63920 34756 63960 34796
rect 78712 34756 78752 34796
rect 78794 34756 78834 34796
rect 78876 34756 78916 34796
rect 78958 34756 78998 34796
rect 79040 34756 79080 34796
rect 93832 34756 93872 34796
rect 93914 34756 93954 34796
rect 93996 34756 94036 34796
rect 94078 34756 94118 34796
rect 94160 34756 94200 34796
rect 4352 34000 4392 34040
rect 4434 34000 4474 34040
rect 4516 34000 4556 34040
rect 4598 34000 4638 34040
rect 4680 34000 4720 34040
rect 19472 34000 19512 34040
rect 19554 34000 19594 34040
rect 19636 34000 19676 34040
rect 19718 34000 19758 34040
rect 19800 34000 19840 34040
rect 34592 34000 34632 34040
rect 34674 34000 34714 34040
rect 34756 34000 34796 34040
rect 34838 34000 34878 34040
rect 34920 34000 34960 34040
rect 49712 34000 49752 34040
rect 49794 34000 49834 34040
rect 49876 34000 49916 34040
rect 49958 34000 49998 34040
rect 50040 34000 50080 34040
rect 64832 34000 64872 34040
rect 64914 34000 64954 34040
rect 64996 34000 65036 34040
rect 65078 34000 65118 34040
rect 65160 34000 65200 34040
rect 79952 34000 79992 34040
rect 80034 34000 80074 34040
rect 80116 34000 80156 34040
rect 80198 34000 80238 34040
rect 80280 34000 80320 34040
rect 95072 34000 95112 34040
rect 95154 34000 95194 34040
rect 95236 34000 95276 34040
rect 95318 34000 95358 34040
rect 95400 34000 95440 34040
rect 3112 33244 3152 33284
rect 3194 33244 3234 33284
rect 3276 33244 3316 33284
rect 3358 33244 3398 33284
rect 3440 33244 3480 33284
rect 18232 33244 18272 33284
rect 18314 33244 18354 33284
rect 18396 33244 18436 33284
rect 18478 33244 18518 33284
rect 18560 33244 18600 33284
rect 33352 33244 33392 33284
rect 33434 33244 33474 33284
rect 33516 33244 33556 33284
rect 33598 33244 33638 33284
rect 33680 33244 33720 33284
rect 48472 33244 48512 33284
rect 48554 33244 48594 33284
rect 48636 33244 48676 33284
rect 48718 33244 48758 33284
rect 48800 33244 48840 33284
rect 63592 33244 63632 33284
rect 63674 33244 63714 33284
rect 63756 33244 63796 33284
rect 63838 33244 63878 33284
rect 63920 33244 63960 33284
rect 78712 33244 78752 33284
rect 78794 33244 78834 33284
rect 78876 33244 78916 33284
rect 78958 33244 78998 33284
rect 79040 33244 79080 33284
rect 93832 33244 93872 33284
rect 93914 33244 93954 33284
rect 93996 33244 94036 33284
rect 94078 33244 94118 33284
rect 94160 33244 94200 33284
rect 4352 32488 4392 32528
rect 4434 32488 4474 32528
rect 4516 32488 4556 32528
rect 4598 32488 4638 32528
rect 4680 32488 4720 32528
rect 19472 32488 19512 32528
rect 19554 32488 19594 32528
rect 19636 32488 19676 32528
rect 19718 32488 19758 32528
rect 19800 32488 19840 32528
rect 34592 32488 34632 32528
rect 34674 32488 34714 32528
rect 34756 32488 34796 32528
rect 34838 32488 34878 32528
rect 34920 32488 34960 32528
rect 49712 32488 49752 32528
rect 49794 32488 49834 32528
rect 49876 32488 49916 32528
rect 49958 32488 49998 32528
rect 50040 32488 50080 32528
rect 64832 32488 64872 32528
rect 64914 32488 64954 32528
rect 64996 32488 65036 32528
rect 65078 32488 65118 32528
rect 65160 32488 65200 32528
rect 79952 32488 79992 32528
rect 80034 32488 80074 32528
rect 80116 32488 80156 32528
rect 80198 32488 80238 32528
rect 80280 32488 80320 32528
rect 95072 32488 95112 32528
rect 95154 32488 95194 32528
rect 95236 32488 95276 32528
rect 95318 32488 95358 32528
rect 95400 32488 95440 32528
rect 3112 31732 3152 31772
rect 3194 31732 3234 31772
rect 3276 31732 3316 31772
rect 3358 31732 3398 31772
rect 3440 31732 3480 31772
rect 18232 31732 18272 31772
rect 18314 31732 18354 31772
rect 18396 31732 18436 31772
rect 18478 31732 18518 31772
rect 18560 31732 18600 31772
rect 33352 31732 33392 31772
rect 33434 31732 33474 31772
rect 33516 31732 33556 31772
rect 33598 31732 33638 31772
rect 33680 31732 33720 31772
rect 48472 31732 48512 31772
rect 48554 31732 48594 31772
rect 48636 31732 48676 31772
rect 48718 31732 48758 31772
rect 48800 31732 48840 31772
rect 63592 31732 63632 31772
rect 63674 31732 63714 31772
rect 63756 31732 63796 31772
rect 63838 31732 63878 31772
rect 63920 31732 63960 31772
rect 78712 31732 78752 31772
rect 78794 31732 78834 31772
rect 78876 31732 78916 31772
rect 78958 31732 78998 31772
rect 79040 31732 79080 31772
rect 93832 31732 93872 31772
rect 93914 31732 93954 31772
rect 93996 31732 94036 31772
rect 94078 31732 94118 31772
rect 94160 31732 94200 31772
rect 4352 30976 4392 31016
rect 4434 30976 4474 31016
rect 4516 30976 4556 31016
rect 4598 30976 4638 31016
rect 4680 30976 4720 31016
rect 19472 30976 19512 31016
rect 19554 30976 19594 31016
rect 19636 30976 19676 31016
rect 19718 30976 19758 31016
rect 19800 30976 19840 31016
rect 34592 30976 34632 31016
rect 34674 30976 34714 31016
rect 34756 30976 34796 31016
rect 34838 30976 34878 31016
rect 34920 30976 34960 31016
rect 49712 30976 49752 31016
rect 49794 30976 49834 31016
rect 49876 30976 49916 31016
rect 49958 30976 49998 31016
rect 50040 30976 50080 31016
rect 64832 30976 64872 31016
rect 64914 30976 64954 31016
rect 64996 30976 65036 31016
rect 65078 30976 65118 31016
rect 65160 30976 65200 31016
rect 79952 30976 79992 31016
rect 80034 30976 80074 31016
rect 80116 30976 80156 31016
rect 80198 30976 80238 31016
rect 80280 30976 80320 31016
rect 95072 30976 95112 31016
rect 95154 30976 95194 31016
rect 95236 30976 95276 31016
rect 95318 30976 95358 31016
rect 95400 30976 95440 31016
rect 3112 30220 3152 30260
rect 3194 30220 3234 30260
rect 3276 30220 3316 30260
rect 3358 30220 3398 30260
rect 3440 30220 3480 30260
rect 18232 30220 18272 30260
rect 18314 30220 18354 30260
rect 18396 30220 18436 30260
rect 18478 30220 18518 30260
rect 18560 30220 18600 30260
rect 33352 30220 33392 30260
rect 33434 30220 33474 30260
rect 33516 30220 33556 30260
rect 33598 30220 33638 30260
rect 33680 30220 33720 30260
rect 48472 30220 48512 30260
rect 48554 30220 48594 30260
rect 48636 30220 48676 30260
rect 48718 30220 48758 30260
rect 48800 30220 48840 30260
rect 63592 30220 63632 30260
rect 63674 30220 63714 30260
rect 63756 30220 63796 30260
rect 63838 30220 63878 30260
rect 63920 30220 63960 30260
rect 78712 30220 78752 30260
rect 78794 30220 78834 30260
rect 78876 30220 78916 30260
rect 78958 30220 78998 30260
rect 79040 30220 79080 30260
rect 93832 30220 93872 30260
rect 93914 30220 93954 30260
rect 93996 30220 94036 30260
rect 94078 30220 94118 30260
rect 94160 30220 94200 30260
rect 4352 29464 4392 29504
rect 4434 29464 4474 29504
rect 4516 29464 4556 29504
rect 4598 29464 4638 29504
rect 4680 29464 4720 29504
rect 19472 29464 19512 29504
rect 19554 29464 19594 29504
rect 19636 29464 19676 29504
rect 19718 29464 19758 29504
rect 19800 29464 19840 29504
rect 34592 29464 34632 29504
rect 34674 29464 34714 29504
rect 34756 29464 34796 29504
rect 34838 29464 34878 29504
rect 34920 29464 34960 29504
rect 49712 29464 49752 29504
rect 49794 29464 49834 29504
rect 49876 29464 49916 29504
rect 49958 29464 49998 29504
rect 50040 29464 50080 29504
rect 64832 29464 64872 29504
rect 64914 29464 64954 29504
rect 64996 29464 65036 29504
rect 65078 29464 65118 29504
rect 65160 29464 65200 29504
rect 79952 29464 79992 29504
rect 80034 29464 80074 29504
rect 80116 29464 80156 29504
rect 80198 29464 80238 29504
rect 80280 29464 80320 29504
rect 95072 29464 95112 29504
rect 95154 29464 95194 29504
rect 95236 29464 95276 29504
rect 95318 29464 95358 29504
rect 95400 29464 95440 29504
rect 3112 28708 3152 28748
rect 3194 28708 3234 28748
rect 3276 28708 3316 28748
rect 3358 28708 3398 28748
rect 3440 28708 3480 28748
rect 18232 28708 18272 28748
rect 18314 28708 18354 28748
rect 18396 28708 18436 28748
rect 18478 28708 18518 28748
rect 18560 28708 18600 28748
rect 33352 28708 33392 28748
rect 33434 28708 33474 28748
rect 33516 28708 33556 28748
rect 33598 28708 33638 28748
rect 33680 28708 33720 28748
rect 48472 28708 48512 28748
rect 48554 28708 48594 28748
rect 48636 28708 48676 28748
rect 48718 28708 48758 28748
rect 48800 28708 48840 28748
rect 63592 28708 63632 28748
rect 63674 28708 63714 28748
rect 63756 28708 63796 28748
rect 63838 28708 63878 28748
rect 63920 28708 63960 28748
rect 78712 28708 78752 28748
rect 78794 28708 78834 28748
rect 78876 28708 78916 28748
rect 78958 28708 78998 28748
rect 79040 28708 79080 28748
rect 93832 28708 93872 28748
rect 93914 28708 93954 28748
rect 93996 28708 94036 28748
rect 94078 28708 94118 28748
rect 94160 28708 94200 28748
rect 4352 27952 4392 27992
rect 4434 27952 4474 27992
rect 4516 27952 4556 27992
rect 4598 27952 4638 27992
rect 4680 27952 4720 27992
rect 19472 27952 19512 27992
rect 19554 27952 19594 27992
rect 19636 27952 19676 27992
rect 19718 27952 19758 27992
rect 19800 27952 19840 27992
rect 34592 27952 34632 27992
rect 34674 27952 34714 27992
rect 34756 27952 34796 27992
rect 34838 27952 34878 27992
rect 34920 27952 34960 27992
rect 49712 27952 49752 27992
rect 49794 27952 49834 27992
rect 49876 27952 49916 27992
rect 49958 27952 49998 27992
rect 50040 27952 50080 27992
rect 64832 27952 64872 27992
rect 64914 27952 64954 27992
rect 64996 27952 65036 27992
rect 65078 27952 65118 27992
rect 65160 27952 65200 27992
rect 79952 27952 79992 27992
rect 80034 27952 80074 27992
rect 80116 27952 80156 27992
rect 80198 27952 80238 27992
rect 80280 27952 80320 27992
rect 95072 27952 95112 27992
rect 95154 27952 95194 27992
rect 95236 27952 95276 27992
rect 95318 27952 95358 27992
rect 95400 27952 95440 27992
rect 3112 27196 3152 27236
rect 3194 27196 3234 27236
rect 3276 27196 3316 27236
rect 3358 27196 3398 27236
rect 3440 27196 3480 27236
rect 18232 27196 18272 27236
rect 18314 27196 18354 27236
rect 18396 27196 18436 27236
rect 18478 27196 18518 27236
rect 18560 27196 18600 27236
rect 33352 27196 33392 27236
rect 33434 27196 33474 27236
rect 33516 27196 33556 27236
rect 33598 27196 33638 27236
rect 33680 27196 33720 27236
rect 48472 27196 48512 27236
rect 48554 27196 48594 27236
rect 48636 27196 48676 27236
rect 48718 27196 48758 27236
rect 48800 27196 48840 27236
rect 63592 27196 63632 27236
rect 63674 27196 63714 27236
rect 63756 27196 63796 27236
rect 63838 27196 63878 27236
rect 63920 27196 63960 27236
rect 78712 27196 78752 27236
rect 78794 27196 78834 27236
rect 78876 27196 78916 27236
rect 78958 27196 78998 27236
rect 79040 27196 79080 27236
rect 93832 27196 93872 27236
rect 93914 27196 93954 27236
rect 93996 27196 94036 27236
rect 94078 27196 94118 27236
rect 94160 27196 94200 27236
rect 4352 26440 4392 26480
rect 4434 26440 4474 26480
rect 4516 26440 4556 26480
rect 4598 26440 4638 26480
rect 4680 26440 4720 26480
rect 19472 26440 19512 26480
rect 19554 26440 19594 26480
rect 19636 26440 19676 26480
rect 19718 26440 19758 26480
rect 19800 26440 19840 26480
rect 34592 26440 34632 26480
rect 34674 26440 34714 26480
rect 34756 26440 34796 26480
rect 34838 26440 34878 26480
rect 34920 26440 34960 26480
rect 49712 26440 49752 26480
rect 49794 26440 49834 26480
rect 49876 26440 49916 26480
rect 49958 26440 49998 26480
rect 50040 26440 50080 26480
rect 64832 26440 64872 26480
rect 64914 26440 64954 26480
rect 64996 26440 65036 26480
rect 65078 26440 65118 26480
rect 65160 26440 65200 26480
rect 79952 26440 79992 26480
rect 80034 26440 80074 26480
rect 80116 26440 80156 26480
rect 80198 26440 80238 26480
rect 80280 26440 80320 26480
rect 95072 26440 95112 26480
rect 95154 26440 95194 26480
rect 95236 26440 95276 26480
rect 95318 26440 95358 26480
rect 95400 26440 95440 26480
rect 3112 25684 3152 25724
rect 3194 25684 3234 25724
rect 3276 25684 3316 25724
rect 3358 25684 3398 25724
rect 3440 25684 3480 25724
rect 18232 25684 18272 25724
rect 18314 25684 18354 25724
rect 18396 25684 18436 25724
rect 18478 25684 18518 25724
rect 18560 25684 18600 25724
rect 33352 25684 33392 25724
rect 33434 25684 33474 25724
rect 33516 25684 33556 25724
rect 33598 25684 33638 25724
rect 33680 25684 33720 25724
rect 48472 25684 48512 25724
rect 48554 25684 48594 25724
rect 48636 25684 48676 25724
rect 48718 25684 48758 25724
rect 48800 25684 48840 25724
rect 63592 25684 63632 25724
rect 63674 25684 63714 25724
rect 63756 25684 63796 25724
rect 63838 25684 63878 25724
rect 63920 25684 63960 25724
rect 78712 25684 78752 25724
rect 78794 25684 78834 25724
rect 78876 25684 78916 25724
rect 78958 25684 78998 25724
rect 79040 25684 79080 25724
rect 93832 25684 93872 25724
rect 93914 25684 93954 25724
rect 93996 25684 94036 25724
rect 94078 25684 94118 25724
rect 94160 25684 94200 25724
rect 4352 24928 4392 24968
rect 4434 24928 4474 24968
rect 4516 24928 4556 24968
rect 4598 24928 4638 24968
rect 4680 24928 4720 24968
rect 19472 24928 19512 24968
rect 19554 24928 19594 24968
rect 19636 24928 19676 24968
rect 19718 24928 19758 24968
rect 19800 24928 19840 24968
rect 34592 24928 34632 24968
rect 34674 24928 34714 24968
rect 34756 24928 34796 24968
rect 34838 24928 34878 24968
rect 34920 24928 34960 24968
rect 49712 24928 49752 24968
rect 49794 24928 49834 24968
rect 49876 24928 49916 24968
rect 49958 24928 49998 24968
rect 50040 24928 50080 24968
rect 64832 24928 64872 24968
rect 64914 24928 64954 24968
rect 64996 24928 65036 24968
rect 65078 24928 65118 24968
rect 65160 24928 65200 24968
rect 79952 24928 79992 24968
rect 80034 24928 80074 24968
rect 80116 24928 80156 24968
rect 80198 24928 80238 24968
rect 80280 24928 80320 24968
rect 95072 24928 95112 24968
rect 95154 24928 95194 24968
rect 95236 24928 95276 24968
rect 95318 24928 95358 24968
rect 95400 24928 95440 24968
rect 3112 24172 3152 24212
rect 3194 24172 3234 24212
rect 3276 24172 3316 24212
rect 3358 24172 3398 24212
rect 3440 24172 3480 24212
rect 18232 24172 18272 24212
rect 18314 24172 18354 24212
rect 18396 24172 18436 24212
rect 18478 24172 18518 24212
rect 18560 24172 18600 24212
rect 33352 24172 33392 24212
rect 33434 24172 33474 24212
rect 33516 24172 33556 24212
rect 33598 24172 33638 24212
rect 33680 24172 33720 24212
rect 48472 24172 48512 24212
rect 48554 24172 48594 24212
rect 48636 24172 48676 24212
rect 48718 24172 48758 24212
rect 48800 24172 48840 24212
rect 63592 24172 63632 24212
rect 63674 24172 63714 24212
rect 63756 24172 63796 24212
rect 63838 24172 63878 24212
rect 63920 24172 63960 24212
rect 78712 24172 78752 24212
rect 78794 24172 78834 24212
rect 78876 24172 78916 24212
rect 78958 24172 78998 24212
rect 79040 24172 79080 24212
rect 93832 24172 93872 24212
rect 93914 24172 93954 24212
rect 93996 24172 94036 24212
rect 94078 24172 94118 24212
rect 94160 24172 94200 24212
rect 4352 23416 4392 23456
rect 4434 23416 4474 23456
rect 4516 23416 4556 23456
rect 4598 23416 4638 23456
rect 4680 23416 4720 23456
rect 19472 23416 19512 23456
rect 19554 23416 19594 23456
rect 19636 23416 19676 23456
rect 19718 23416 19758 23456
rect 19800 23416 19840 23456
rect 34592 23416 34632 23456
rect 34674 23416 34714 23456
rect 34756 23416 34796 23456
rect 34838 23416 34878 23456
rect 34920 23416 34960 23456
rect 49712 23416 49752 23456
rect 49794 23416 49834 23456
rect 49876 23416 49916 23456
rect 49958 23416 49998 23456
rect 50040 23416 50080 23456
rect 64832 23416 64872 23456
rect 64914 23416 64954 23456
rect 64996 23416 65036 23456
rect 65078 23416 65118 23456
rect 65160 23416 65200 23456
rect 79952 23416 79992 23456
rect 80034 23416 80074 23456
rect 80116 23416 80156 23456
rect 80198 23416 80238 23456
rect 80280 23416 80320 23456
rect 95072 23416 95112 23456
rect 95154 23416 95194 23456
rect 95236 23416 95276 23456
rect 95318 23416 95358 23456
rect 95400 23416 95440 23456
rect 3112 22660 3152 22700
rect 3194 22660 3234 22700
rect 3276 22660 3316 22700
rect 3358 22660 3398 22700
rect 3440 22660 3480 22700
rect 18232 22660 18272 22700
rect 18314 22660 18354 22700
rect 18396 22660 18436 22700
rect 18478 22660 18518 22700
rect 18560 22660 18600 22700
rect 33352 22660 33392 22700
rect 33434 22660 33474 22700
rect 33516 22660 33556 22700
rect 33598 22660 33638 22700
rect 33680 22660 33720 22700
rect 48472 22660 48512 22700
rect 48554 22660 48594 22700
rect 48636 22660 48676 22700
rect 48718 22660 48758 22700
rect 48800 22660 48840 22700
rect 63592 22660 63632 22700
rect 63674 22660 63714 22700
rect 63756 22660 63796 22700
rect 63838 22660 63878 22700
rect 63920 22660 63960 22700
rect 78712 22660 78752 22700
rect 78794 22660 78834 22700
rect 78876 22660 78916 22700
rect 78958 22660 78998 22700
rect 79040 22660 79080 22700
rect 93832 22660 93872 22700
rect 93914 22660 93954 22700
rect 93996 22660 94036 22700
rect 94078 22660 94118 22700
rect 94160 22660 94200 22700
rect 4352 21904 4392 21944
rect 4434 21904 4474 21944
rect 4516 21904 4556 21944
rect 4598 21904 4638 21944
rect 4680 21904 4720 21944
rect 19472 21904 19512 21944
rect 19554 21904 19594 21944
rect 19636 21904 19676 21944
rect 19718 21904 19758 21944
rect 19800 21904 19840 21944
rect 34592 21904 34632 21944
rect 34674 21904 34714 21944
rect 34756 21904 34796 21944
rect 34838 21904 34878 21944
rect 34920 21904 34960 21944
rect 49712 21904 49752 21944
rect 49794 21904 49834 21944
rect 49876 21904 49916 21944
rect 49958 21904 49998 21944
rect 50040 21904 50080 21944
rect 64832 21904 64872 21944
rect 64914 21904 64954 21944
rect 64996 21904 65036 21944
rect 65078 21904 65118 21944
rect 65160 21904 65200 21944
rect 79952 21904 79992 21944
rect 80034 21904 80074 21944
rect 80116 21904 80156 21944
rect 80198 21904 80238 21944
rect 80280 21904 80320 21944
rect 95072 21904 95112 21944
rect 95154 21904 95194 21944
rect 95236 21904 95276 21944
rect 95318 21904 95358 21944
rect 95400 21904 95440 21944
rect 3112 21148 3152 21188
rect 3194 21148 3234 21188
rect 3276 21148 3316 21188
rect 3358 21148 3398 21188
rect 3440 21148 3480 21188
rect 18232 21148 18272 21188
rect 18314 21148 18354 21188
rect 18396 21148 18436 21188
rect 18478 21148 18518 21188
rect 18560 21148 18600 21188
rect 33352 21148 33392 21188
rect 33434 21148 33474 21188
rect 33516 21148 33556 21188
rect 33598 21148 33638 21188
rect 33680 21148 33720 21188
rect 48472 21148 48512 21188
rect 48554 21148 48594 21188
rect 48636 21148 48676 21188
rect 48718 21148 48758 21188
rect 48800 21148 48840 21188
rect 63592 21148 63632 21188
rect 63674 21148 63714 21188
rect 63756 21148 63796 21188
rect 63838 21148 63878 21188
rect 63920 21148 63960 21188
rect 78712 21148 78752 21188
rect 78794 21148 78834 21188
rect 78876 21148 78916 21188
rect 78958 21148 78998 21188
rect 79040 21148 79080 21188
rect 93832 21148 93872 21188
rect 93914 21148 93954 21188
rect 93996 21148 94036 21188
rect 94078 21148 94118 21188
rect 94160 21148 94200 21188
rect 4352 20392 4392 20432
rect 4434 20392 4474 20432
rect 4516 20392 4556 20432
rect 4598 20392 4638 20432
rect 4680 20392 4720 20432
rect 19472 20392 19512 20432
rect 19554 20392 19594 20432
rect 19636 20392 19676 20432
rect 19718 20392 19758 20432
rect 19800 20392 19840 20432
rect 34592 20392 34632 20432
rect 34674 20392 34714 20432
rect 34756 20392 34796 20432
rect 34838 20392 34878 20432
rect 34920 20392 34960 20432
rect 49712 20392 49752 20432
rect 49794 20392 49834 20432
rect 49876 20392 49916 20432
rect 49958 20392 49998 20432
rect 50040 20392 50080 20432
rect 64832 20392 64872 20432
rect 64914 20392 64954 20432
rect 64996 20392 65036 20432
rect 65078 20392 65118 20432
rect 65160 20392 65200 20432
rect 79952 20392 79992 20432
rect 80034 20392 80074 20432
rect 80116 20392 80156 20432
rect 80198 20392 80238 20432
rect 80280 20392 80320 20432
rect 95072 20392 95112 20432
rect 95154 20392 95194 20432
rect 95236 20392 95276 20432
rect 95318 20392 95358 20432
rect 95400 20392 95440 20432
rect 3112 19636 3152 19676
rect 3194 19636 3234 19676
rect 3276 19636 3316 19676
rect 3358 19636 3398 19676
rect 3440 19636 3480 19676
rect 18232 19636 18272 19676
rect 18314 19636 18354 19676
rect 18396 19636 18436 19676
rect 18478 19636 18518 19676
rect 18560 19636 18600 19676
rect 33352 19636 33392 19676
rect 33434 19636 33474 19676
rect 33516 19636 33556 19676
rect 33598 19636 33638 19676
rect 33680 19636 33720 19676
rect 48472 19636 48512 19676
rect 48554 19636 48594 19676
rect 48636 19636 48676 19676
rect 48718 19636 48758 19676
rect 48800 19636 48840 19676
rect 63592 19636 63632 19676
rect 63674 19636 63714 19676
rect 63756 19636 63796 19676
rect 63838 19636 63878 19676
rect 63920 19636 63960 19676
rect 78712 19636 78752 19676
rect 78794 19636 78834 19676
rect 78876 19636 78916 19676
rect 78958 19636 78998 19676
rect 79040 19636 79080 19676
rect 93832 19636 93872 19676
rect 93914 19636 93954 19676
rect 93996 19636 94036 19676
rect 94078 19636 94118 19676
rect 94160 19636 94200 19676
rect 4352 18880 4392 18920
rect 4434 18880 4474 18920
rect 4516 18880 4556 18920
rect 4598 18880 4638 18920
rect 4680 18880 4720 18920
rect 19472 18880 19512 18920
rect 19554 18880 19594 18920
rect 19636 18880 19676 18920
rect 19718 18880 19758 18920
rect 19800 18880 19840 18920
rect 34592 18880 34632 18920
rect 34674 18880 34714 18920
rect 34756 18880 34796 18920
rect 34838 18880 34878 18920
rect 34920 18880 34960 18920
rect 49712 18880 49752 18920
rect 49794 18880 49834 18920
rect 49876 18880 49916 18920
rect 49958 18880 49998 18920
rect 50040 18880 50080 18920
rect 64832 18880 64872 18920
rect 64914 18880 64954 18920
rect 64996 18880 65036 18920
rect 65078 18880 65118 18920
rect 65160 18880 65200 18920
rect 79952 18880 79992 18920
rect 80034 18880 80074 18920
rect 80116 18880 80156 18920
rect 80198 18880 80238 18920
rect 80280 18880 80320 18920
rect 95072 18880 95112 18920
rect 95154 18880 95194 18920
rect 95236 18880 95276 18920
rect 95318 18880 95358 18920
rect 95400 18880 95440 18920
rect 3112 18124 3152 18164
rect 3194 18124 3234 18164
rect 3276 18124 3316 18164
rect 3358 18124 3398 18164
rect 3440 18124 3480 18164
rect 18232 18124 18272 18164
rect 18314 18124 18354 18164
rect 18396 18124 18436 18164
rect 18478 18124 18518 18164
rect 18560 18124 18600 18164
rect 33352 18124 33392 18164
rect 33434 18124 33474 18164
rect 33516 18124 33556 18164
rect 33598 18124 33638 18164
rect 33680 18124 33720 18164
rect 48472 18124 48512 18164
rect 48554 18124 48594 18164
rect 48636 18124 48676 18164
rect 48718 18124 48758 18164
rect 48800 18124 48840 18164
rect 63592 18124 63632 18164
rect 63674 18124 63714 18164
rect 63756 18124 63796 18164
rect 63838 18124 63878 18164
rect 63920 18124 63960 18164
rect 78712 18124 78752 18164
rect 78794 18124 78834 18164
rect 78876 18124 78916 18164
rect 78958 18124 78998 18164
rect 79040 18124 79080 18164
rect 93832 18124 93872 18164
rect 93914 18124 93954 18164
rect 93996 18124 94036 18164
rect 94078 18124 94118 18164
rect 94160 18124 94200 18164
rect 4352 17368 4392 17408
rect 4434 17368 4474 17408
rect 4516 17368 4556 17408
rect 4598 17368 4638 17408
rect 4680 17368 4720 17408
rect 19472 17368 19512 17408
rect 19554 17368 19594 17408
rect 19636 17368 19676 17408
rect 19718 17368 19758 17408
rect 19800 17368 19840 17408
rect 34592 17368 34632 17408
rect 34674 17368 34714 17408
rect 34756 17368 34796 17408
rect 34838 17368 34878 17408
rect 34920 17368 34960 17408
rect 49712 17368 49752 17408
rect 49794 17368 49834 17408
rect 49876 17368 49916 17408
rect 49958 17368 49998 17408
rect 50040 17368 50080 17408
rect 64832 17368 64872 17408
rect 64914 17368 64954 17408
rect 64996 17368 65036 17408
rect 65078 17368 65118 17408
rect 65160 17368 65200 17408
rect 79952 17368 79992 17408
rect 80034 17368 80074 17408
rect 80116 17368 80156 17408
rect 80198 17368 80238 17408
rect 80280 17368 80320 17408
rect 95072 17368 95112 17408
rect 95154 17368 95194 17408
rect 95236 17368 95276 17408
rect 95318 17368 95358 17408
rect 95400 17368 95440 17408
rect 3112 16612 3152 16652
rect 3194 16612 3234 16652
rect 3276 16612 3316 16652
rect 3358 16612 3398 16652
rect 3440 16612 3480 16652
rect 18232 16612 18272 16652
rect 18314 16612 18354 16652
rect 18396 16612 18436 16652
rect 18478 16612 18518 16652
rect 18560 16612 18600 16652
rect 33352 16612 33392 16652
rect 33434 16612 33474 16652
rect 33516 16612 33556 16652
rect 33598 16612 33638 16652
rect 33680 16612 33720 16652
rect 48472 16612 48512 16652
rect 48554 16612 48594 16652
rect 48636 16612 48676 16652
rect 48718 16612 48758 16652
rect 48800 16612 48840 16652
rect 63592 16612 63632 16652
rect 63674 16612 63714 16652
rect 63756 16612 63796 16652
rect 63838 16612 63878 16652
rect 63920 16612 63960 16652
rect 78712 16612 78752 16652
rect 78794 16612 78834 16652
rect 78876 16612 78916 16652
rect 78958 16612 78998 16652
rect 79040 16612 79080 16652
rect 93832 16612 93872 16652
rect 93914 16612 93954 16652
rect 93996 16612 94036 16652
rect 94078 16612 94118 16652
rect 94160 16612 94200 16652
rect 4352 15856 4392 15896
rect 4434 15856 4474 15896
rect 4516 15856 4556 15896
rect 4598 15856 4638 15896
rect 4680 15856 4720 15896
rect 19472 15856 19512 15896
rect 19554 15856 19594 15896
rect 19636 15856 19676 15896
rect 19718 15856 19758 15896
rect 19800 15856 19840 15896
rect 34592 15856 34632 15896
rect 34674 15856 34714 15896
rect 34756 15856 34796 15896
rect 34838 15856 34878 15896
rect 34920 15856 34960 15896
rect 49712 15856 49752 15896
rect 49794 15856 49834 15896
rect 49876 15856 49916 15896
rect 49958 15856 49998 15896
rect 50040 15856 50080 15896
rect 64832 15856 64872 15896
rect 64914 15856 64954 15896
rect 64996 15856 65036 15896
rect 65078 15856 65118 15896
rect 65160 15856 65200 15896
rect 79952 15856 79992 15896
rect 80034 15856 80074 15896
rect 80116 15856 80156 15896
rect 80198 15856 80238 15896
rect 80280 15856 80320 15896
rect 95072 15856 95112 15896
rect 95154 15856 95194 15896
rect 95236 15856 95276 15896
rect 95318 15856 95358 15896
rect 95400 15856 95440 15896
rect 3112 15100 3152 15140
rect 3194 15100 3234 15140
rect 3276 15100 3316 15140
rect 3358 15100 3398 15140
rect 3440 15100 3480 15140
rect 18232 15100 18272 15140
rect 18314 15100 18354 15140
rect 18396 15100 18436 15140
rect 18478 15100 18518 15140
rect 18560 15100 18600 15140
rect 33352 15100 33392 15140
rect 33434 15100 33474 15140
rect 33516 15100 33556 15140
rect 33598 15100 33638 15140
rect 33680 15100 33720 15140
rect 48472 15100 48512 15140
rect 48554 15100 48594 15140
rect 48636 15100 48676 15140
rect 48718 15100 48758 15140
rect 48800 15100 48840 15140
rect 63592 15100 63632 15140
rect 63674 15100 63714 15140
rect 63756 15100 63796 15140
rect 63838 15100 63878 15140
rect 63920 15100 63960 15140
rect 78712 15100 78752 15140
rect 78794 15100 78834 15140
rect 78876 15100 78916 15140
rect 78958 15100 78998 15140
rect 79040 15100 79080 15140
rect 93832 15100 93872 15140
rect 93914 15100 93954 15140
rect 93996 15100 94036 15140
rect 94078 15100 94118 15140
rect 94160 15100 94200 15140
rect 4352 14344 4392 14384
rect 4434 14344 4474 14384
rect 4516 14344 4556 14384
rect 4598 14344 4638 14384
rect 4680 14344 4720 14384
rect 19472 14344 19512 14384
rect 19554 14344 19594 14384
rect 19636 14344 19676 14384
rect 19718 14344 19758 14384
rect 19800 14344 19840 14384
rect 34592 14344 34632 14384
rect 34674 14344 34714 14384
rect 34756 14344 34796 14384
rect 34838 14344 34878 14384
rect 34920 14344 34960 14384
rect 49712 14344 49752 14384
rect 49794 14344 49834 14384
rect 49876 14344 49916 14384
rect 49958 14344 49998 14384
rect 50040 14344 50080 14384
rect 64832 14344 64872 14384
rect 64914 14344 64954 14384
rect 64996 14344 65036 14384
rect 65078 14344 65118 14384
rect 65160 14344 65200 14384
rect 79952 14344 79992 14384
rect 80034 14344 80074 14384
rect 80116 14344 80156 14384
rect 80198 14344 80238 14384
rect 80280 14344 80320 14384
rect 95072 14344 95112 14384
rect 95154 14344 95194 14384
rect 95236 14344 95276 14384
rect 95318 14344 95358 14384
rect 95400 14344 95440 14384
rect 3112 13588 3152 13628
rect 3194 13588 3234 13628
rect 3276 13588 3316 13628
rect 3358 13588 3398 13628
rect 3440 13588 3480 13628
rect 18232 13588 18272 13628
rect 18314 13588 18354 13628
rect 18396 13588 18436 13628
rect 18478 13588 18518 13628
rect 18560 13588 18600 13628
rect 33352 13588 33392 13628
rect 33434 13588 33474 13628
rect 33516 13588 33556 13628
rect 33598 13588 33638 13628
rect 33680 13588 33720 13628
rect 48472 13588 48512 13628
rect 48554 13588 48594 13628
rect 48636 13588 48676 13628
rect 48718 13588 48758 13628
rect 48800 13588 48840 13628
rect 63592 13588 63632 13628
rect 63674 13588 63714 13628
rect 63756 13588 63796 13628
rect 63838 13588 63878 13628
rect 63920 13588 63960 13628
rect 78712 13588 78752 13628
rect 78794 13588 78834 13628
rect 78876 13588 78916 13628
rect 78958 13588 78998 13628
rect 79040 13588 79080 13628
rect 93832 13588 93872 13628
rect 93914 13588 93954 13628
rect 93996 13588 94036 13628
rect 94078 13588 94118 13628
rect 94160 13588 94200 13628
rect 4352 12832 4392 12872
rect 4434 12832 4474 12872
rect 4516 12832 4556 12872
rect 4598 12832 4638 12872
rect 4680 12832 4720 12872
rect 19472 12832 19512 12872
rect 19554 12832 19594 12872
rect 19636 12832 19676 12872
rect 19718 12832 19758 12872
rect 19800 12832 19840 12872
rect 34592 12832 34632 12872
rect 34674 12832 34714 12872
rect 34756 12832 34796 12872
rect 34838 12832 34878 12872
rect 34920 12832 34960 12872
rect 49712 12832 49752 12872
rect 49794 12832 49834 12872
rect 49876 12832 49916 12872
rect 49958 12832 49998 12872
rect 50040 12832 50080 12872
rect 64832 12832 64872 12872
rect 64914 12832 64954 12872
rect 64996 12832 65036 12872
rect 65078 12832 65118 12872
rect 65160 12832 65200 12872
rect 79952 12832 79992 12872
rect 80034 12832 80074 12872
rect 80116 12832 80156 12872
rect 80198 12832 80238 12872
rect 80280 12832 80320 12872
rect 95072 12832 95112 12872
rect 95154 12832 95194 12872
rect 95236 12832 95276 12872
rect 95318 12832 95358 12872
rect 95400 12832 95440 12872
rect 3112 12076 3152 12116
rect 3194 12076 3234 12116
rect 3276 12076 3316 12116
rect 3358 12076 3398 12116
rect 3440 12076 3480 12116
rect 18232 12076 18272 12116
rect 18314 12076 18354 12116
rect 18396 12076 18436 12116
rect 18478 12076 18518 12116
rect 18560 12076 18600 12116
rect 33352 12076 33392 12116
rect 33434 12076 33474 12116
rect 33516 12076 33556 12116
rect 33598 12076 33638 12116
rect 33680 12076 33720 12116
rect 48472 12076 48512 12116
rect 48554 12076 48594 12116
rect 48636 12076 48676 12116
rect 48718 12076 48758 12116
rect 48800 12076 48840 12116
rect 63592 12076 63632 12116
rect 63674 12076 63714 12116
rect 63756 12076 63796 12116
rect 63838 12076 63878 12116
rect 63920 12076 63960 12116
rect 78712 12076 78752 12116
rect 78794 12076 78834 12116
rect 78876 12076 78916 12116
rect 78958 12076 78998 12116
rect 79040 12076 79080 12116
rect 93832 12076 93872 12116
rect 93914 12076 93954 12116
rect 93996 12076 94036 12116
rect 94078 12076 94118 12116
rect 94160 12076 94200 12116
rect 4352 11320 4392 11360
rect 4434 11320 4474 11360
rect 4516 11320 4556 11360
rect 4598 11320 4638 11360
rect 4680 11320 4720 11360
rect 19472 11320 19512 11360
rect 19554 11320 19594 11360
rect 19636 11320 19676 11360
rect 19718 11320 19758 11360
rect 19800 11320 19840 11360
rect 34592 11320 34632 11360
rect 34674 11320 34714 11360
rect 34756 11320 34796 11360
rect 34838 11320 34878 11360
rect 34920 11320 34960 11360
rect 49712 11320 49752 11360
rect 49794 11320 49834 11360
rect 49876 11320 49916 11360
rect 49958 11320 49998 11360
rect 50040 11320 50080 11360
rect 64832 11320 64872 11360
rect 64914 11320 64954 11360
rect 64996 11320 65036 11360
rect 65078 11320 65118 11360
rect 65160 11320 65200 11360
rect 79952 11320 79992 11360
rect 80034 11320 80074 11360
rect 80116 11320 80156 11360
rect 80198 11320 80238 11360
rect 80280 11320 80320 11360
rect 95072 11320 95112 11360
rect 95154 11320 95194 11360
rect 95236 11320 95276 11360
rect 95318 11320 95358 11360
rect 95400 11320 95440 11360
rect 3112 10564 3152 10604
rect 3194 10564 3234 10604
rect 3276 10564 3316 10604
rect 3358 10564 3398 10604
rect 3440 10564 3480 10604
rect 18232 10564 18272 10604
rect 18314 10564 18354 10604
rect 18396 10564 18436 10604
rect 18478 10564 18518 10604
rect 18560 10564 18600 10604
rect 33352 10564 33392 10604
rect 33434 10564 33474 10604
rect 33516 10564 33556 10604
rect 33598 10564 33638 10604
rect 33680 10564 33720 10604
rect 48472 10564 48512 10604
rect 48554 10564 48594 10604
rect 48636 10564 48676 10604
rect 48718 10564 48758 10604
rect 48800 10564 48840 10604
rect 63592 10564 63632 10604
rect 63674 10564 63714 10604
rect 63756 10564 63796 10604
rect 63838 10564 63878 10604
rect 63920 10564 63960 10604
rect 78712 10564 78752 10604
rect 78794 10564 78834 10604
rect 78876 10564 78916 10604
rect 78958 10564 78998 10604
rect 79040 10564 79080 10604
rect 93832 10564 93872 10604
rect 93914 10564 93954 10604
rect 93996 10564 94036 10604
rect 94078 10564 94118 10604
rect 94160 10564 94200 10604
rect 4352 9808 4392 9848
rect 4434 9808 4474 9848
rect 4516 9808 4556 9848
rect 4598 9808 4638 9848
rect 4680 9808 4720 9848
rect 19472 9808 19512 9848
rect 19554 9808 19594 9848
rect 19636 9808 19676 9848
rect 19718 9808 19758 9848
rect 19800 9808 19840 9848
rect 34592 9808 34632 9848
rect 34674 9808 34714 9848
rect 34756 9808 34796 9848
rect 34838 9808 34878 9848
rect 34920 9808 34960 9848
rect 49712 9808 49752 9848
rect 49794 9808 49834 9848
rect 49876 9808 49916 9848
rect 49958 9808 49998 9848
rect 50040 9808 50080 9848
rect 64832 9808 64872 9848
rect 64914 9808 64954 9848
rect 64996 9808 65036 9848
rect 65078 9808 65118 9848
rect 65160 9808 65200 9848
rect 79952 9808 79992 9848
rect 80034 9808 80074 9848
rect 80116 9808 80156 9848
rect 80198 9808 80238 9848
rect 80280 9808 80320 9848
rect 95072 9808 95112 9848
rect 95154 9808 95194 9848
rect 95236 9808 95276 9848
rect 95318 9808 95358 9848
rect 95400 9808 95440 9848
rect 3112 9052 3152 9092
rect 3194 9052 3234 9092
rect 3276 9052 3316 9092
rect 3358 9052 3398 9092
rect 3440 9052 3480 9092
rect 18232 9052 18272 9092
rect 18314 9052 18354 9092
rect 18396 9052 18436 9092
rect 18478 9052 18518 9092
rect 18560 9052 18600 9092
rect 33352 9052 33392 9092
rect 33434 9052 33474 9092
rect 33516 9052 33556 9092
rect 33598 9052 33638 9092
rect 33680 9052 33720 9092
rect 48472 9052 48512 9092
rect 48554 9052 48594 9092
rect 48636 9052 48676 9092
rect 48718 9052 48758 9092
rect 48800 9052 48840 9092
rect 63592 9052 63632 9092
rect 63674 9052 63714 9092
rect 63756 9052 63796 9092
rect 63838 9052 63878 9092
rect 63920 9052 63960 9092
rect 78712 9052 78752 9092
rect 78794 9052 78834 9092
rect 78876 9052 78916 9092
rect 78958 9052 78998 9092
rect 79040 9052 79080 9092
rect 93832 9052 93872 9092
rect 93914 9052 93954 9092
rect 93996 9052 94036 9092
rect 94078 9052 94118 9092
rect 94160 9052 94200 9092
rect 4352 8296 4392 8336
rect 4434 8296 4474 8336
rect 4516 8296 4556 8336
rect 4598 8296 4638 8336
rect 4680 8296 4720 8336
rect 19472 8296 19512 8336
rect 19554 8296 19594 8336
rect 19636 8296 19676 8336
rect 19718 8296 19758 8336
rect 19800 8296 19840 8336
rect 34592 8296 34632 8336
rect 34674 8296 34714 8336
rect 34756 8296 34796 8336
rect 34838 8296 34878 8336
rect 34920 8296 34960 8336
rect 49712 8296 49752 8336
rect 49794 8296 49834 8336
rect 49876 8296 49916 8336
rect 49958 8296 49998 8336
rect 50040 8296 50080 8336
rect 64832 8296 64872 8336
rect 64914 8296 64954 8336
rect 64996 8296 65036 8336
rect 65078 8296 65118 8336
rect 65160 8296 65200 8336
rect 79952 8296 79992 8336
rect 80034 8296 80074 8336
rect 80116 8296 80156 8336
rect 80198 8296 80238 8336
rect 80280 8296 80320 8336
rect 95072 8296 95112 8336
rect 95154 8296 95194 8336
rect 95236 8296 95276 8336
rect 95318 8296 95358 8336
rect 95400 8296 95440 8336
rect 3112 7540 3152 7580
rect 3194 7540 3234 7580
rect 3276 7540 3316 7580
rect 3358 7540 3398 7580
rect 3440 7540 3480 7580
rect 18232 7540 18272 7580
rect 18314 7540 18354 7580
rect 18396 7540 18436 7580
rect 18478 7540 18518 7580
rect 18560 7540 18600 7580
rect 33352 7540 33392 7580
rect 33434 7540 33474 7580
rect 33516 7540 33556 7580
rect 33598 7540 33638 7580
rect 33680 7540 33720 7580
rect 48472 7540 48512 7580
rect 48554 7540 48594 7580
rect 48636 7540 48676 7580
rect 48718 7540 48758 7580
rect 48800 7540 48840 7580
rect 63592 7540 63632 7580
rect 63674 7540 63714 7580
rect 63756 7540 63796 7580
rect 63838 7540 63878 7580
rect 63920 7540 63960 7580
rect 78712 7540 78752 7580
rect 78794 7540 78834 7580
rect 78876 7540 78916 7580
rect 78958 7540 78998 7580
rect 79040 7540 79080 7580
rect 93832 7540 93872 7580
rect 93914 7540 93954 7580
rect 93996 7540 94036 7580
rect 94078 7540 94118 7580
rect 94160 7540 94200 7580
rect 4352 6784 4392 6824
rect 4434 6784 4474 6824
rect 4516 6784 4556 6824
rect 4598 6784 4638 6824
rect 4680 6784 4720 6824
rect 19472 6784 19512 6824
rect 19554 6784 19594 6824
rect 19636 6784 19676 6824
rect 19718 6784 19758 6824
rect 19800 6784 19840 6824
rect 34592 6784 34632 6824
rect 34674 6784 34714 6824
rect 34756 6784 34796 6824
rect 34838 6784 34878 6824
rect 34920 6784 34960 6824
rect 49712 6784 49752 6824
rect 49794 6784 49834 6824
rect 49876 6784 49916 6824
rect 49958 6784 49998 6824
rect 50040 6784 50080 6824
rect 64832 6784 64872 6824
rect 64914 6784 64954 6824
rect 64996 6784 65036 6824
rect 65078 6784 65118 6824
rect 65160 6784 65200 6824
rect 79952 6784 79992 6824
rect 80034 6784 80074 6824
rect 80116 6784 80156 6824
rect 80198 6784 80238 6824
rect 80280 6784 80320 6824
rect 95072 6784 95112 6824
rect 95154 6784 95194 6824
rect 95236 6784 95276 6824
rect 95318 6784 95358 6824
rect 95400 6784 95440 6824
rect 3112 6028 3152 6068
rect 3194 6028 3234 6068
rect 3276 6028 3316 6068
rect 3358 6028 3398 6068
rect 3440 6028 3480 6068
rect 18232 6028 18272 6068
rect 18314 6028 18354 6068
rect 18396 6028 18436 6068
rect 18478 6028 18518 6068
rect 18560 6028 18600 6068
rect 33352 6028 33392 6068
rect 33434 6028 33474 6068
rect 33516 6028 33556 6068
rect 33598 6028 33638 6068
rect 33680 6028 33720 6068
rect 48472 6028 48512 6068
rect 48554 6028 48594 6068
rect 48636 6028 48676 6068
rect 48718 6028 48758 6068
rect 48800 6028 48840 6068
rect 63592 6028 63632 6068
rect 63674 6028 63714 6068
rect 63756 6028 63796 6068
rect 63838 6028 63878 6068
rect 63920 6028 63960 6068
rect 78712 6028 78752 6068
rect 78794 6028 78834 6068
rect 78876 6028 78916 6068
rect 78958 6028 78998 6068
rect 79040 6028 79080 6068
rect 93832 6028 93872 6068
rect 93914 6028 93954 6068
rect 93996 6028 94036 6068
rect 94078 6028 94118 6068
rect 94160 6028 94200 6068
rect 4352 5272 4392 5312
rect 4434 5272 4474 5312
rect 4516 5272 4556 5312
rect 4598 5272 4638 5312
rect 4680 5272 4720 5312
rect 19472 5272 19512 5312
rect 19554 5272 19594 5312
rect 19636 5272 19676 5312
rect 19718 5272 19758 5312
rect 19800 5272 19840 5312
rect 34592 5272 34632 5312
rect 34674 5272 34714 5312
rect 34756 5272 34796 5312
rect 34838 5272 34878 5312
rect 34920 5272 34960 5312
rect 49712 5272 49752 5312
rect 49794 5272 49834 5312
rect 49876 5272 49916 5312
rect 49958 5272 49998 5312
rect 50040 5272 50080 5312
rect 64832 5272 64872 5312
rect 64914 5272 64954 5312
rect 64996 5272 65036 5312
rect 65078 5272 65118 5312
rect 65160 5272 65200 5312
rect 79952 5272 79992 5312
rect 80034 5272 80074 5312
rect 80116 5272 80156 5312
rect 80198 5272 80238 5312
rect 80280 5272 80320 5312
rect 95072 5272 95112 5312
rect 95154 5272 95194 5312
rect 95236 5272 95276 5312
rect 95318 5272 95358 5312
rect 95400 5272 95440 5312
rect 3112 4516 3152 4556
rect 3194 4516 3234 4556
rect 3276 4516 3316 4556
rect 3358 4516 3398 4556
rect 3440 4516 3480 4556
rect 18232 4516 18272 4556
rect 18314 4516 18354 4556
rect 18396 4516 18436 4556
rect 18478 4516 18518 4556
rect 18560 4516 18600 4556
rect 33352 4516 33392 4556
rect 33434 4516 33474 4556
rect 33516 4516 33556 4556
rect 33598 4516 33638 4556
rect 33680 4516 33720 4556
rect 48472 4516 48512 4556
rect 48554 4516 48594 4556
rect 48636 4516 48676 4556
rect 48718 4516 48758 4556
rect 48800 4516 48840 4556
rect 63592 4516 63632 4556
rect 63674 4516 63714 4556
rect 63756 4516 63796 4556
rect 63838 4516 63878 4556
rect 63920 4516 63960 4556
rect 78712 4516 78752 4556
rect 78794 4516 78834 4556
rect 78876 4516 78916 4556
rect 78958 4516 78998 4556
rect 79040 4516 79080 4556
rect 93832 4516 93872 4556
rect 93914 4516 93954 4556
rect 93996 4516 94036 4556
rect 94078 4516 94118 4556
rect 94160 4516 94200 4556
rect 4352 3760 4392 3800
rect 4434 3760 4474 3800
rect 4516 3760 4556 3800
rect 4598 3760 4638 3800
rect 4680 3760 4720 3800
rect 19472 3760 19512 3800
rect 19554 3760 19594 3800
rect 19636 3760 19676 3800
rect 19718 3760 19758 3800
rect 19800 3760 19840 3800
rect 34592 3760 34632 3800
rect 34674 3760 34714 3800
rect 34756 3760 34796 3800
rect 34838 3760 34878 3800
rect 34920 3760 34960 3800
rect 49712 3760 49752 3800
rect 49794 3760 49834 3800
rect 49876 3760 49916 3800
rect 49958 3760 49998 3800
rect 50040 3760 50080 3800
rect 64832 3760 64872 3800
rect 64914 3760 64954 3800
rect 64996 3760 65036 3800
rect 65078 3760 65118 3800
rect 65160 3760 65200 3800
rect 79952 3760 79992 3800
rect 80034 3760 80074 3800
rect 80116 3760 80156 3800
rect 80198 3760 80238 3800
rect 80280 3760 80320 3800
rect 95072 3760 95112 3800
rect 95154 3760 95194 3800
rect 95236 3760 95276 3800
rect 95318 3760 95358 3800
rect 95400 3760 95440 3800
rect 3112 3004 3152 3044
rect 3194 3004 3234 3044
rect 3276 3004 3316 3044
rect 3358 3004 3398 3044
rect 3440 3004 3480 3044
rect 18232 3004 18272 3044
rect 18314 3004 18354 3044
rect 18396 3004 18436 3044
rect 18478 3004 18518 3044
rect 18560 3004 18600 3044
rect 33352 3004 33392 3044
rect 33434 3004 33474 3044
rect 33516 3004 33556 3044
rect 33598 3004 33638 3044
rect 33680 3004 33720 3044
rect 48472 3004 48512 3044
rect 48554 3004 48594 3044
rect 48636 3004 48676 3044
rect 48718 3004 48758 3044
rect 48800 3004 48840 3044
rect 63592 3004 63632 3044
rect 63674 3004 63714 3044
rect 63756 3004 63796 3044
rect 63838 3004 63878 3044
rect 63920 3004 63960 3044
rect 78712 3004 78752 3044
rect 78794 3004 78834 3044
rect 78876 3004 78916 3044
rect 78958 3004 78998 3044
rect 79040 3004 79080 3044
rect 93832 3004 93872 3044
rect 93914 3004 93954 3044
rect 93996 3004 94036 3044
rect 94078 3004 94118 3044
rect 94160 3004 94200 3044
rect 4352 2248 4392 2288
rect 4434 2248 4474 2288
rect 4516 2248 4556 2288
rect 4598 2248 4638 2288
rect 4680 2248 4720 2288
rect 19472 2248 19512 2288
rect 19554 2248 19594 2288
rect 19636 2248 19676 2288
rect 19718 2248 19758 2288
rect 19800 2248 19840 2288
rect 34592 2248 34632 2288
rect 34674 2248 34714 2288
rect 34756 2248 34796 2288
rect 34838 2248 34878 2288
rect 34920 2248 34960 2288
rect 49712 2248 49752 2288
rect 49794 2248 49834 2288
rect 49876 2248 49916 2288
rect 49958 2248 49998 2288
rect 50040 2248 50080 2288
rect 64832 2248 64872 2288
rect 64914 2248 64954 2288
rect 64996 2248 65036 2288
rect 65078 2248 65118 2288
rect 65160 2248 65200 2288
rect 79952 2248 79992 2288
rect 80034 2248 80074 2288
rect 80116 2248 80156 2288
rect 80198 2248 80238 2288
rect 80280 2248 80320 2288
rect 95072 2248 95112 2288
rect 95154 2248 95194 2288
rect 95236 2248 95276 2288
rect 95318 2248 95358 2288
rect 95400 2248 95440 2288
rect 3112 1492 3152 1532
rect 3194 1492 3234 1532
rect 3276 1492 3316 1532
rect 3358 1492 3398 1532
rect 3440 1492 3480 1532
rect 18232 1492 18272 1532
rect 18314 1492 18354 1532
rect 18396 1492 18436 1532
rect 18478 1492 18518 1532
rect 18560 1492 18600 1532
rect 33352 1492 33392 1532
rect 33434 1492 33474 1532
rect 33516 1492 33556 1532
rect 33598 1492 33638 1532
rect 33680 1492 33720 1532
rect 48472 1492 48512 1532
rect 48554 1492 48594 1532
rect 48636 1492 48676 1532
rect 48718 1492 48758 1532
rect 48800 1492 48840 1532
rect 63592 1492 63632 1532
rect 63674 1492 63714 1532
rect 63756 1492 63796 1532
rect 63838 1492 63878 1532
rect 63920 1492 63960 1532
rect 78712 1492 78752 1532
rect 78794 1492 78834 1532
rect 78876 1492 78916 1532
rect 78958 1492 78998 1532
rect 79040 1492 79080 1532
rect 93832 1492 93872 1532
rect 93914 1492 93954 1532
rect 93996 1492 94036 1532
rect 94078 1492 94118 1532
rect 94160 1492 94200 1532
rect 4352 736 4392 776
rect 4434 736 4474 776
rect 4516 736 4556 776
rect 4598 736 4638 776
rect 4680 736 4720 776
rect 19472 736 19512 776
rect 19554 736 19594 776
rect 19636 736 19676 776
rect 19718 736 19758 776
rect 19800 736 19840 776
rect 34592 736 34632 776
rect 34674 736 34714 776
rect 34756 736 34796 776
rect 34838 736 34878 776
rect 34920 736 34960 776
rect 49712 736 49752 776
rect 49794 736 49834 776
rect 49876 736 49916 776
rect 49958 736 49998 776
rect 50040 736 50080 776
rect 64832 736 64872 776
rect 64914 736 64954 776
rect 64996 736 65036 776
rect 65078 736 65118 776
rect 65160 736 65200 776
rect 79952 736 79992 776
rect 80034 736 80074 776
rect 80116 736 80156 776
rect 80198 736 80238 776
rect 80280 736 80320 776
rect 95072 736 95112 776
rect 95154 736 95194 776
rect 95236 736 95276 776
rect 95318 736 95358 776
rect 95400 736 95440 776
<< metal4 >>
rect 4352 38576 4720 38585
rect 4392 38536 4434 38576
rect 4474 38536 4516 38576
rect 4556 38536 4598 38576
rect 4638 38536 4680 38576
rect 4352 38527 4720 38536
rect 19472 38576 19840 38585
rect 19512 38536 19554 38576
rect 19594 38536 19636 38576
rect 19676 38536 19718 38576
rect 19758 38536 19800 38576
rect 19472 38527 19840 38536
rect 34592 38576 34960 38585
rect 34632 38536 34674 38576
rect 34714 38536 34756 38576
rect 34796 38536 34838 38576
rect 34878 38536 34920 38576
rect 34592 38527 34960 38536
rect 49712 38576 50080 38585
rect 49752 38536 49794 38576
rect 49834 38536 49876 38576
rect 49916 38536 49958 38576
rect 49998 38536 50040 38576
rect 49712 38527 50080 38536
rect 64832 38576 65200 38585
rect 64872 38536 64914 38576
rect 64954 38536 64996 38576
rect 65036 38536 65078 38576
rect 65118 38536 65160 38576
rect 64832 38527 65200 38536
rect 79952 38576 80320 38585
rect 79992 38536 80034 38576
rect 80074 38536 80116 38576
rect 80156 38536 80198 38576
rect 80238 38536 80280 38576
rect 79952 38527 80320 38536
rect 95072 38576 95440 38585
rect 95112 38536 95154 38576
rect 95194 38536 95236 38576
rect 95276 38536 95318 38576
rect 95358 38536 95400 38576
rect 95072 38527 95440 38536
rect 3112 37820 3480 37829
rect 3152 37780 3194 37820
rect 3234 37780 3276 37820
rect 3316 37780 3358 37820
rect 3398 37780 3440 37820
rect 3112 37771 3480 37780
rect 18232 37820 18600 37829
rect 18272 37780 18314 37820
rect 18354 37780 18396 37820
rect 18436 37780 18478 37820
rect 18518 37780 18560 37820
rect 18232 37771 18600 37780
rect 33352 37820 33720 37829
rect 33392 37780 33434 37820
rect 33474 37780 33516 37820
rect 33556 37780 33598 37820
rect 33638 37780 33680 37820
rect 33352 37771 33720 37780
rect 48472 37820 48840 37829
rect 48512 37780 48554 37820
rect 48594 37780 48636 37820
rect 48676 37780 48718 37820
rect 48758 37780 48800 37820
rect 48472 37771 48840 37780
rect 63592 37820 63960 37829
rect 63632 37780 63674 37820
rect 63714 37780 63756 37820
rect 63796 37780 63838 37820
rect 63878 37780 63920 37820
rect 63592 37771 63960 37780
rect 78712 37820 79080 37829
rect 78752 37780 78794 37820
rect 78834 37780 78876 37820
rect 78916 37780 78958 37820
rect 78998 37780 79040 37820
rect 78712 37771 79080 37780
rect 93832 37820 94200 37829
rect 93872 37780 93914 37820
rect 93954 37780 93996 37820
rect 94036 37780 94078 37820
rect 94118 37780 94160 37820
rect 93832 37771 94200 37780
rect 4352 37064 4720 37073
rect 4392 37024 4434 37064
rect 4474 37024 4516 37064
rect 4556 37024 4598 37064
rect 4638 37024 4680 37064
rect 4352 37015 4720 37024
rect 19472 37064 19840 37073
rect 19512 37024 19554 37064
rect 19594 37024 19636 37064
rect 19676 37024 19718 37064
rect 19758 37024 19800 37064
rect 19472 37015 19840 37024
rect 34592 37064 34960 37073
rect 34632 37024 34674 37064
rect 34714 37024 34756 37064
rect 34796 37024 34838 37064
rect 34878 37024 34920 37064
rect 34592 37015 34960 37024
rect 49712 37064 50080 37073
rect 49752 37024 49794 37064
rect 49834 37024 49876 37064
rect 49916 37024 49958 37064
rect 49998 37024 50040 37064
rect 49712 37015 50080 37024
rect 64832 37064 65200 37073
rect 64872 37024 64914 37064
rect 64954 37024 64996 37064
rect 65036 37024 65078 37064
rect 65118 37024 65160 37064
rect 64832 37015 65200 37024
rect 79952 37064 80320 37073
rect 79992 37024 80034 37064
rect 80074 37024 80116 37064
rect 80156 37024 80198 37064
rect 80238 37024 80280 37064
rect 79952 37015 80320 37024
rect 95072 37064 95440 37073
rect 95112 37024 95154 37064
rect 95194 37024 95236 37064
rect 95276 37024 95318 37064
rect 95358 37024 95400 37064
rect 95072 37015 95440 37024
rect 3112 36308 3480 36317
rect 3152 36268 3194 36308
rect 3234 36268 3276 36308
rect 3316 36268 3358 36308
rect 3398 36268 3440 36308
rect 3112 36259 3480 36268
rect 18232 36308 18600 36317
rect 18272 36268 18314 36308
rect 18354 36268 18396 36308
rect 18436 36268 18478 36308
rect 18518 36268 18560 36308
rect 18232 36259 18600 36268
rect 33352 36308 33720 36317
rect 33392 36268 33434 36308
rect 33474 36268 33516 36308
rect 33556 36268 33598 36308
rect 33638 36268 33680 36308
rect 33352 36259 33720 36268
rect 48472 36308 48840 36317
rect 48512 36268 48554 36308
rect 48594 36268 48636 36308
rect 48676 36268 48718 36308
rect 48758 36268 48800 36308
rect 48472 36259 48840 36268
rect 63592 36308 63960 36317
rect 63632 36268 63674 36308
rect 63714 36268 63756 36308
rect 63796 36268 63838 36308
rect 63878 36268 63920 36308
rect 63592 36259 63960 36268
rect 78712 36308 79080 36317
rect 78752 36268 78794 36308
rect 78834 36268 78876 36308
rect 78916 36268 78958 36308
rect 78998 36268 79040 36308
rect 78712 36259 79080 36268
rect 93832 36308 94200 36317
rect 93872 36268 93914 36308
rect 93954 36268 93996 36308
rect 94036 36268 94078 36308
rect 94118 36268 94160 36308
rect 93832 36259 94200 36268
rect 4352 35552 4720 35561
rect 4392 35512 4434 35552
rect 4474 35512 4516 35552
rect 4556 35512 4598 35552
rect 4638 35512 4680 35552
rect 4352 35503 4720 35512
rect 19472 35552 19840 35561
rect 19512 35512 19554 35552
rect 19594 35512 19636 35552
rect 19676 35512 19718 35552
rect 19758 35512 19800 35552
rect 19472 35503 19840 35512
rect 34592 35552 34960 35561
rect 34632 35512 34674 35552
rect 34714 35512 34756 35552
rect 34796 35512 34838 35552
rect 34878 35512 34920 35552
rect 34592 35503 34960 35512
rect 49712 35552 50080 35561
rect 49752 35512 49794 35552
rect 49834 35512 49876 35552
rect 49916 35512 49958 35552
rect 49998 35512 50040 35552
rect 49712 35503 50080 35512
rect 64832 35552 65200 35561
rect 64872 35512 64914 35552
rect 64954 35512 64996 35552
rect 65036 35512 65078 35552
rect 65118 35512 65160 35552
rect 64832 35503 65200 35512
rect 79952 35552 80320 35561
rect 79992 35512 80034 35552
rect 80074 35512 80116 35552
rect 80156 35512 80198 35552
rect 80238 35512 80280 35552
rect 79952 35503 80320 35512
rect 95072 35552 95440 35561
rect 95112 35512 95154 35552
rect 95194 35512 95236 35552
rect 95276 35512 95318 35552
rect 95358 35512 95400 35552
rect 95072 35503 95440 35512
rect 3112 34796 3480 34805
rect 3152 34756 3194 34796
rect 3234 34756 3276 34796
rect 3316 34756 3358 34796
rect 3398 34756 3440 34796
rect 3112 34747 3480 34756
rect 18232 34796 18600 34805
rect 18272 34756 18314 34796
rect 18354 34756 18396 34796
rect 18436 34756 18478 34796
rect 18518 34756 18560 34796
rect 18232 34747 18600 34756
rect 33352 34796 33720 34805
rect 33392 34756 33434 34796
rect 33474 34756 33516 34796
rect 33556 34756 33598 34796
rect 33638 34756 33680 34796
rect 33352 34747 33720 34756
rect 48472 34796 48840 34805
rect 48512 34756 48554 34796
rect 48594 34756 48636 34796
rect 48676 34756 48718 34796
rect 48758 34756 48800 34796
rect 48472 34747 48840 34756
rect 63592 34796 63960 34805
rect 63632 34756 63674 34796
rect 63714 34756 63756 34796
rect 63796 34756 63838 34796
rect 63878 34756 63920 34796
rect 63592 34747 63960 34756
rect 78712 34796 79080 34805
rect 78752 34756 78794 34796
rect 78834 34756 78876 34796
rect 78916 34756 78958 34796
rect 78998 34756 79040 34796
rect 78712 34747 79080 34756
rect 93832 34796 94200 34805
rect 93872 34756 93914 34796
rect 93954 34756 93996 34796
rect 94036 34756 94078 34796
rect 94118 34756 94160 34796
rect 93832 34747 94200 34756
rect 4352 34040 4720 34049
rect 4392 34000 4434 34040
rect 4474 34000 4516 34040
rect 4556 34000 4598 34040
rect 4638 34000 4680 34040
rect 4352 33991 4720 34000
rect 19472 34040 19840 34049
rect 19512 34000 19554 34040
rect 19594 34000 19636 34040
rect 19676 34000 19718 34040
rect 19758 34000 19800 34040
rect 19472 33991 19840 34000
rect 34592 34040 34960 34049
rect 34632 34000 34674 34040
rect 34714 34000 34756 34040
rect 34796 34000 34838 34040
rect 34878 34000 34920 34040
rect 34592 33991 34960 34000
rect 49712 34040 50080 34049
rect 49752 34000 49794 34040
rect 49834 34000 49876 34040
rect 49916 34000 49958 34040
rect 49998 34000 50040 34040
rect 49712 33991 50080 34000
rect 64832 34040 65200 34049
rect 64872 34000 64914 34040
rect 64954 34000 64996 34040
rect 65036 34000 65078 34040
rect 65118 34000 65160 34040
rect 64832 33991 65200 34000
rect 79952 34040 80320 34049
rect 79992 34000 80034 34040
rect 80074 34000 80116 34040
rect 80156 34000 80198 34040
rect 80238 34000 80280 34040
rect 79952 33991 80320 34000
rect 95072 34040 95440 34049
rect 95112 34000 95154 34040
rect 95194 34000 95236 34040
rect 95276 34000 95318 34040
rect 95358 34000 95400 34040
rect 95072 33991 95440 34000
rect 3112 33284 3480 33293
rect 3152 33244 3194 33284
rect 3234 33244 3276 33284
rect 3316 33244 3358 33284
rect 3398 33244 3440 33284
rect 3112 33235 3480 33244
rect 18232 33284 18600 33293
rect 18272 33244 18314 33284
rect 18354 33244 18396 33284
rect 18436 33244 18478 33284
rect 18518 33244 18560 33284
rect 18232 33235 18600 33244
rect 33352 33284 33720 33293
rect 33392 33244 33434 33284
rect 33474 33244 33516 33284
rect 33556 33244 33598 33284
rect 33638 33244 33680 33284
rect 33352 33235 33720 33244
rect 48472 33284 48840 33293
rect 48512 33244 48554 33284
rect 48594 33244 48636 33284
rect 48676 33244 48718 33284
rect 48758 33244 48800 33284
rect 48472 33235 48840 33244
rect 63592 33284 63960 33293
rect 63632 33244 63674 33284
rect 63714 33244 63756 33284
rect 63796 33244 63838 33284
rect 63878 33244 63920 33284
rect 63592 33235 63960 33244
rect 78712 33284 79080 33293
rect 78752 33244 78794 33284
rect 78834 33244 78876 33284
rect 78916 33244 78958 33284
rect 78998 33244 79040 33284
rect 78712 33235 79080 33244
rect 93832 33284 94200 33293
rect 93872 33244 93914 33284
rect 93954 33244 93996 33284
rect 94036 33244 94078 33284
rect 94118 33244 94160 33284
rect 93832 33235 94200 33244
rect 4352 32528 4720 32537
rect 4392 32488 4434 32528
rect 4474 32488 4516 32528
rect 4556 32488 4598 32528
rect 4638 32488 4680 32528
rect 4352 32479 4720 32488
rect 19472 32528 19840 32537
rect 19512 32488 19554 32528
rect 19594 32488 19636 32528
rect 19676 32488 19718 32528
rect 19758 32488 19800 32528
rect 19472 32479 19840 32488
rect 34592 32528 34960 32537
rect 34632 32488 34674 32528
rect 34714 32488 34756 32528
rect 34796 32488 34838 32528
rect 34878 32488 34920 32528
rect 34592 32479 34960 32488
rect 49712 32528 50080 32537
rect 49752 32488 49794 32528
rect 49834 32488 49876 32528
rect 49916 32488 49958 32528
rect 49998 32488 50040 32528
rect 49712 32479 50080 32488
rect 64832 32528 65200 32537
rect 64872 32488 64914 32528
rect 64954 32488 64996 32528
rect 65036 32488 65078 32528
rect 65118 32488 65160 32528
rect 64832 32479 65200 32488
rect 79952 32528 80320 32537
rect 79992 32488 80034 32528
rect 80074 32488 80116 32528
rect 80156 32488 80198 32528
rect 80238 32488 80280 32528
rect 79952 32479 80320 32488
rect 95072 32528 95440 32537
rect 95112 32488 95154 32528
rect 95194 32488 95236 32528
rect 95276 32488 95318 32528
rect 95358 32488 95400 32528
rect 95072 32479 95440 32488
rect 3112 31772 3480 31781
rect 3152 31732 3194 31772
rect 3234 31732 3276 31772
rect 3316 31732 3358 31772
rect 3398 31732 3440 31772
rect 3112 31723 3480 31732
rect 18232 31772 18600 31781
rect 18272 31732 18314 31772
rect 18354 31732 18396 31772
rect 18436 31732 18478 31772
rect 18518 31732 18560 31772
rect 18232 31723 18600 31732
rect 33352 31772 33720 31781
rect 33392 31732 33434 31772
rect 33474 31732 33516 31772
rect 33556 31732 33598 31772
rect 33638 31732 33680 31772
rect 33352 31723 33720 31732
rect 48472 31772 48840 31781
rect 48512 31732 48554 31772
rect 48594 31732 48636 31772
rect 48676 31732 48718 31772
rect 48758 31732 48800 31772
rect 48472 31723 48840 31732
rect 63592 31772 63960 31781
rect 63632 31732 63674 31772
rect 63714 31732 63756 31772
rect 63796 31732 63838 31772
rect 63878 31732 63920 31772
rect 63592 31723 63960 31732
rect 78712 31772 79080 31781
rect 78752 31732 78794 31772
rect 78834 31732 78876 31772
rect 78916 31732 78958 31772
rect 78998 31732 79040 31772
rect 78712 31723 79080 31732
rect 93832 31772 94200 31781
rect 93872 31732 93914 31772
rect 93954 31732 93996 31772
rect 94036 31732 94078 31772
rect 94118 31732 94160 31772
rect 93832 31723 94200 31732
rect 4352 31016 4720 31025
rect 4392 30976 4434 31016
rect 4474 30976 4516 31016
rect 4556 30976 4598 31016
rect 4638 30976 4680 31016
rect 4352 30967 4720 30976
rect 19472 31016 19840 31025
rect 19512 30976 19554 31016
rect 19594 30976 19636 31016
rect 19676 30976 19718 31016
rect 19758 30976 19800 31016
rect 19472 30967 19840 30976
rect 34592 31016 34960 31025
rect 34632 30976 34674 31016
rect 34714 30976 34756 31016
rect 34796 30976 34838 31016
rect 34878 30976 34920 31016
rect 34592 30967 34960 30976
rect 49712 31016 50080 31025
rect 49752 30976 49794 31016
rect 49834 30976 49876 31016
rect 49916 30976 49958 31016
rect 49998 30976 50040 31016
rect 49712 30967 50080 30976
rect 64832 31016 65200 31025
rect 64872 30976 64914 31016
rect 64954 30976 64996 31016
rect 65036 30976 65078 31016
rect 65118 30976 65160 31016
rect 64832 30967 65200 30976
rect 79952 31016 80320 31025
rect 79992 30976 80034 31016
rect 80074 30976 80116 31016
rect 80156 30976 80198 31016
rect 80238 30976 80280 31016
rect 79952 30967 80320 30976
rect 95072 31016 95440 31025
rect 95112 30976 95154 31016
rect 95194 30976 95236 31016
rect 95276 30976 95318 31016
rect 95358 30976 95400 31016
rect 95072 30967 95440 30976
rect 3112 30260 3480 30269
rect 3152 30220 3194 30260
rect 3234 30220 3276 30260
rect 3316 30220 3358 30260
rect 3398 30220 3440 30260
rect 3112 30211 3480 30220
rect 18232 30260 18600 30269
rect 18272 30220 18314 30260
rect 18354 30220 18396 30260
rect 18436 30220 18478 30260
rect 18518 30220 18560 30260
rect 18232 30211 18600 30220
rect 33352 30260 33720 30269
rect 33392 30220 33434 30260
rect 33474 30220 33516 30260
rect 33556 30220 33598 30260
rect 33638 30220 33680 30260
rect 33352 30211 33720 30220
rect 48472 30260 48840 30269
rect 48512 30220 48554 30260
rect 48594 30220 48636 30260
rect 48676 30220 48718 30260
rect 48758 30220 48800 30260
rect 48472 30211 48840 30220
rect 63592 30260 63960 30269
rect 63632 30220 63674 30260
rect 63714 30220 63756 30260
rect 63796 30220 63838 30260
rect 63878 30220 63920 30260
rect 63592 30211 63960 30220
rect 78712 30260 79080 30269
rect 78752 30220 78794 30260
rect 78834 30220 78876 30260
rect 78916 30220 78958 30260
rect 78998 30220 79040 30260
rect 78712 30211 79080 30220
rect 93832 30260 94200 30269
rect 93872 30220 93914 30260
rect 93954 30220 93996 30260
rect 94036 30220 94078 30260
rect 94118 30220 94160 30260
rect 93832 30211 94200 30220
rect 4352 29504 4720 29513
rect 4392 29464 4434 29504
rect 4474 29464 4516 29504
rect 4556 29464 4598 29504
rect 4638 29464 4680 29504
rect 4352 29455 4720 29464
rect 19472 29504 19840 29513
rect 19512 29464 19554 29504
rect 19594 29464 19636 29504
rect 19676 29464 19718 29504
rect 19758 29464 19800 29504
rect 19472 29455 19840 29464
rect 34592 29504 34960 29513
rect 34632 29464 34674 29504
rect 34714 29464 34756 29504
rect 34796 29464 34838 29504
rect 34878 29464 34920 29504
rect 34592 29455 34960 29464
rect 49712 29504 50080 29513
rect 49752 29464 49794 29504
rect 49834 29464 49876 29504
rect 49916 29464 49958 29504
rect 49998 29464 50040 29504
rect 49712 29455 50080 29464
rect 64832 29504 65200 29513
rect 64872 29464 64914 29504
rect 64954 29464 64996 29504
rect 65036 29464 65078 29504
rect 65118 29464 65160 29504
rect 64832 29455 65200 29464
rect 79952 29504 80320 29513
rect 79992 29464 80034 29504
rect 80074 29464 80116 29504
rect 80156 29464 80198 29504
rect 80238 29464 80280 29504
rect 79952 29455 80320 29464
rect 95072 29504 95440 29513
rect 95112 29464 95154 29504
rect 95194 29464 95236 29504
rect 95276 29464 95318 29504
rect 95358 29464 95400 29504
rect 95072 29455 95440 29464
rect 3112 28748 3480 28757
rect 3152 28708 3194 28748
rect 3234 28708 3276 28748
rect 3316 28708 3358 28748
rect 3398 28708 3440 28748
rect 3112 28699 3480 28708
rect 18232 28748 18600 28757
rect 18272 28708 18314 28748
rect 18354 28708 18396 28748
rect 18436 28708 18478 28748
rect 18518 28708 18560 28748
rect 18232 28699 18600 28708
rect 33352 28748 33720 28757
rect 33392 28708 33434 28748
rect 33474 28708 33516 28748
rect 33556 28708 33598 28748
rect 33638 28708 33680 28748
rect 33352 28699 33720 28708
rect 48472 28748 48840 28757
rect 48512 28708 48554 28748
rect 48594 28708 48636 28748
rect 48676 28708 48718 28748
rect 48758 28708 48800 28748
rect 48472 28699 48840 28708
rect 63592 28748 63960 28757
rect 63632 28708 63674 28748
rect 63714 28708 63756 28748
rect 63796 28708 63838 28748
rect 63878 28708 63920 28748
rect 63592 28699 63960 28708
rect 78712 28748 79080 28757
rect 78752 28708 78794 28748
rect 78834 28708 78876 28748
rect 78916 28708 78958 28748
rect 78998 28708 79040 28748
rect 78712 28699 79080 28708
rect 93832 28748 94200 28757
rect 93872 28708 93914 28748
rect 93954 28708 93996 28748
rect 94036 28708 94078 28748
rect 94118 28708 94160 28748
rect 93832 28699 94200 28708
rect 4352 27992 4720 28001
rect 4392 27952 4434 27992
rect 4474 27952 4516 27992
rect 4556 27952 4598 27992
rect 4638 27952 4680 27992
rect 4352 27943 4720 27952
rect 19472 27992 19840 28001
rect 19512 27952 19554 27992
rect 19594 27952 19636 27992
rect 19676 27952 19718 27992
rect 19758 27952 19800 27992
rect 19472 27943 19840 27952
rect 34592 27992 34960 28001
rect 34632 27952 34674 27992
rect 34714 27952 34756 27992
rect 34796 27952 34838 27992
rect 34878 27952 34920 27992
rect 34592 27943 34960 27952
rect 49712 27992 50080 28001
rect 49752 27952 49794 27992
rect 49834 27952 49876 27992
rect 49916 27952 49958 27992
rect 49998 27952 50040 27992
rect 49712 27943 50080 27952
rect 64832 27992 65200 28001
rect 64872 27952 64914 27992
rect 64954 27952 64996 27992
rect 65036 27952 65078 27992
rect 65118 27952 65160 27992
rect 64832 27943 65200 27952
rect 79952 27992 80320 28001
rect 79992 27952 80034 27992
rect 80074 27952 80116 27992
rect 80156 27952 80198 27992
rect 80238 27952 80280 27992
rect 79952 27943 80320 27952
rect 95072 27992 95440 28001
rect 95112 27952 95154 27992
rect 95194 27952 95236 27992
rect 95276 27952 95318 27992
rect 95358 27952 95400 27992
rect 95072 27943 95440 27952
rect 3112 27236 3480 27245
rect 3152 27196 3194 27236
rect 3234 27196 3276 27236
rect 3316 27196 3358 27236
rect 3398 27196 3440 27236
rect 3112 27187 3480 27196
rect 18232 27236 18600 27245
rect 18272 27196 18314 27236
rect 18354 27196 18396 27236
rect 18436 27196 18478 27236
rect 18518 27196 18560 27236
rect 18232 27187 18600 27196
rect 33352 27236 33720 27245
rect 33392 27196 33434 27236
rect 33474 27196 33516 27236
rect 33556 27196 33598 27236
rect 33638 27196 33680 27236
rect 33352 27187 33720 27196
rect 48472 27236 48840 27245
rect 48512 27196 48554 27236
rect 48594 27196 48636 27236
rect 48676 27196 48718 27236
rect 48758 27196 48800 27236
rect 48472 27187 48840 27196
rect 63592 27236 63960 27245
rect 63632 27196 63674 27236
rect 63714 27196 63756 27236
rect 63796 27196 63838 27236
rect 63878 27196 63920 27236
rect 63592 27187 63960 27196
rect 78712 27236 79080 27245
rect 78752 27196 78794 27236
rect 78834 27196 78876 27236
rect 78916 27196 78958 27236
rect 78998 27196 79040 27236
rect 78712 27187 79080 27196
rect 93832 27236 94200 27245
rect 93872 27196 93914 27236
rect 93954 27196 93996 27236
rect 94036 27196 94078 27236
rect 94118 27196 94160 27236
rect 93832 27187 94200 27196
rect 4352 26480 4720 26489
rect 4392 26440 4434 26480
rect 4474 26440 4516 26480
rect 4556 26440 4598 26480
rect 4638 26440 4680 26480
rect 4352 26431 4720 26440
rect 19472 26480 19840 26489
rect 19512 26440 19554 26480
rect 19594 26440 19636 26480
rect 19676 26440 19718 26480
rect 19758 26440 19800 26480
rect 19472 26431 19840 26440
rect 34592 26480 34960 26489
rect 34632 26440 34674 26480
rect 34714 26440 34756 26480
rect 34796 26440 34838 26480
rect 34878 26440 34920 26480
rect 34592 26431 34960 26440
rect 49712 26480 50080 26489
rect 49752 26440 49794 26480
rect 49834 26440 49876 26480
rect 49916 26440 49958 26480
rect 49998 26440 50040 26480
rect 49712 26431 50080 26440
rect 64832 26480 65200 26489
rect 64872 26440 64914 26480
rect 64954 26440 64996 26480
rect 65036 26440 65078 26480
rect 65118 26440 65160 26480
rect 64832 26431 65200 26440
rect 79952 26480 80320 26489
rect 79992 26440 80034 26480
rect 80074 26440 80116 26480
rect 80156 26440 80198 26480
rect 80238 26440 80280 26480
rect 79952 26431 80320 26440
rect 95072 26480 95440 26489
rect 95112 26440 95154 26480
rect 95194 26440 95236 26480
rect 95276 26440 95318 26480
rect 95358 26440 95400 26480
rect 95072 26431 95440 26440
rect 3112 25724 3480 25733
rect 3152 25684 3194 25724
rect 3234 25684 3276 25724
rect 3316 25684 3358 25724
rect 3398 25684 3440 25724
rect 3112 25675 3480 25684
rect 18232 25724 18600 25733
rect 18272 25684 18314 25724
rect 18354 25684 18396 25724
rect 18436 25684 18478 25724
rect 18518 25684 18560 25724
rect 18232 25675 18600 25684
rect 33352 25724 33720 25733
rect 33392 25684 33434 25724
rect 33474 25684 33516 25724
rect 33556 25684 33598 25724
rect 33638 25684 33680 25724
rect 33352 25675 33720 25684
rect 48472 25724 48840 25733
rect 48512 25684 48554 25724
rect 48594 25684 48636 25724
rect 48676 25684 48718 25724
rect 48758 25684 48800 25724
rect 48472 25675 48840 25684
rect 63592 25724 63960 25733
rect 63632 25684 63674 25724
rect 63714 25684 63756 25724
rect 63796 25684 63838 25724
rect 63878 25684 63920 25724
rect 63592 25675 63960 25684
rect 78712 25724 79080 25733
rect 78752 25684 78794 25724
rect 78834 25684 78876 25724
rect 78916 25684 78958 25724
rect 78998 25684 79040 25724
rect 78712 25675 79080 25684
rect 93832 25724 94200 25733
rect 93872 25684 93914 25724
rect 93954 25684 93996 25724
rect 94036 25684 94078 25724
rect 94118 25684 94160 25724
rect 93832 25675 94200 25684
rect 4352 24968 4720 24977
rect 4392 24928 4434 24968
rect 4474 24928 4516 24968
rect 4556 24928 4598 24968
rect 4638 24928 4680 24968
rect 4352 24919 4720 24928
rect 19472 24968 19840 24977
rect 19512 24928 19554 24968
rect 19594 24928 19636 24968
rect 19676 24928 19718 24968
rect 19758 24928 19800 24968
rect 19472 24919 19840 24928
rect 34592 24968 34960 24977
rect 34632 24928 34674 24968
rect 34714 24928 34756 24968
rect 34796 24928 34838 24968
rect 34878 24928 34920 24968
rect 34592 24919 34960 24928
rect 49712 24968 50080 24977
rect 49752 24928 49794 24968
rect 49834 24928 49876 24968
rect 49916 24928 49958 24968
rect 49998 24928 50040 24968
rect 49712 24919 50080 24928
rect 64832 24968 65200 24977
rect 64872 24928 64914 24968
rect 64954 24928 64996 24968
rect 65036 24928 65078 24968
rect 65118 24928 65160 24968
rect 64832 24919 65200 24928
rect 79952 24968 80320 24977
rect 79992 24928 80034 24968
rect 80074 24928 80116 24968
rect 80156 24928 80198 24968
rect 80238 24928 80280 24968
rect 79952 24919 80320 24928
rect 95072 24968 95440 24977
rect 95112 24928 95154 24968
rect 95194 24928 95236 24968
rect 95276 24928 95318 24968
rect 95358 24928 95400 24968
rect 95072 24919 95440 24928
rect 3112 24212 3480 24221
rect 3152 24172 3194 24212
rect 3234 24172 3276 24212
rect 3316 24172 3358 24212
rect 3398 24172 3440 24212
rect 3112 24163 3480 24172
rect 18232 24212 18600 24221
rect 18272 24172 18314 24212
rect 18354 24172 18396 24212
rect 18436 24172 18478 24212
rect 18518 24172 18560 24212
rect 18232 24163 18600 24172
rect 33352 24212 33720 24221
rect 33392 24172 33434 24212
rect 33474 24172 33516 24212
rect 33556 24172 33598 24212
rect 33638 24172 33680 24212
rect 33352 24163 33720 24172
rect 48472 24212 48840 24221
rect 48512 24172 48554 24212
rect 48594 24172 48636 24212
rect 48676 24172 48718 24212
rect 48758 24172 48800 24212
rect 48472 24163 48840 24172
rect 63592 24212 63960 24221
rect 63632 24172 63674 24212
rect 63714 24172 63756 24212
rect 63796 24172 63838 24212
rect 63878 24172 63920 24212
rect 63592 24163 63960 24172
rect 78712 24212 79080 24221
rect 78752 24172 78794 24212
rect 78834 24172 78876 24212
rect 78916 24172 78958 24212
rect 78998 24172 79040 24212
rect 78712 24163 79080 24172
rect 93832 24212 94200 24221
rect 93872 24172 93914 24212
rect 93954 24172 93996 24212
rect 94036 24172 94078 24212
rect 94118 24172 94160 24212
rect 93832 24163 94200 24172
rect 4352 23456 4720 23465
rect 4392 23416 4434 23456
rect 4474 23416 4516 23456
rect 4556 23416 4598 23456
rect 4638 23416 4680 23456
rect 4352 23407 4720 23416
rect 19472 23456 19840 23465
rect 19512 23416 19554 23456
rect 19594 23416 19636 23456
rect 19676 23416 19718 23456
rect 19758 23416 19800 23456
rect 19472 23407 19840 23416
rect 34592 23456 34960 23465
rect 34632 23416 34674 23456
rect 34714 23416 34756 23456
rect 34796 23416 34838 23456
rect 34878 23416 34920 23456
rect 34592 23407 34960 23416
rect 49712 23456 50080 23465
rect 49752 23416 49794 23456
rect 49834 23416 49876 23456
rect 49916 23416 49958 23456
rect 49998 23416 50040 23456
rect 49712 23407 50080 23416
rect 64832 23456 65200 23465
rect 64872 23416 64914 23456
rect 64954 23416 64996 23456
rect 65036 23416 65078 23456
rect 65118 23416 65160 23456
rect 64832 23407 65200 23416
rect 79952 23456 80320 23465
rect 79992 23416 80034 23456
rect 80074 23416 80116 23456
rect 80156 23416 80198 23456
rect 80238 23416 80280 23456
rect 79952 23407 80320 23416
rect 95072 23456 95440 23465
rect 95112 23416 95154 23456
rect 95194 23416 95236 23456
rect 95276 23416 95318 23456
rect 95358 23416 95400 23456
rect 95072 23407 95440 23416
rect 3112 22700 3480 22709
rect 3152 22660 3194 22700
rect 3234 22660 3276 22700
rect 3316 22660 3358 22700
rect 3398 22660 3440 22700
rect 3112 22651 3480 22660
rect 18232 22700 18600 22709
rect 18272 22660 18314 22700
rect 18354 22660 18396 22700
rect 18436 22660 18478 22700
rect 18518 22660 18560 22700
rect 18232 22651 18600 22660
rect 33352 22700 33720 22709
rect 33392 22660 33434 22700
rect 33474 22660 33516 22700
rect 33556 22660 33598 22700
rect 33638 22660 33680 22700
rect 33352 22651 33720 22660
rect 48472 22700 48840 22709
rect 48512 22660 48554 22700
rect 48594 22660 48636 22700
rect 48676 22660 48718 22700
rect 48758 22660 48800 22700
rect 48472 22651 48840 22660
rect 63592 22700 63960 22709
rect 63632 22660 63674 22700
rect 63714 22660 63756 22700
rect 63796 22660 63838 22700
rect 63878 22660 63920 22700
rect 63592 22651 63960 22660
rect 78712 22700 79080 22709
rect 78752 22660 78794 22700
rect 78834 22660 78876 22700
rect 78916 22660 78958 22700
rect 78998 22660 79040 22700
rect 78712 22651 79080 22660
rect 93832 22700 94200 22709
rect 93872 22660 93914 22700
rect 93954 22660 93996 22700
rect 94036 22660 94078 22700
rect 94118 22660 94160 22700
rect 93832 22651 94200 22660
rect 4352 21944 4720 21953
rect 4392 21904 4434 21944
rect 4474 21904 4516 21944
rect 4556 21904 4598 21944
rect 4638 21904 4680 21944
rect 4352 21895 4720 21904
rect 19472 21944 19840 21953
rect 19512 21904 19554 21944
rect 19594 21904 19636 21944
rect 19676 21904 19718 21944
rect 19758 21904 19800 21944
rect 19472 21895 19840 21904
rect 34592 21944 34960 21953
rect 34632 21904 34674 21944
rect 34714 21904 34756 21944
rect 34796 21904 34838 21944
rect 34878 21904 34920 21944
rect 34592 21895 34960 21904
rect 49712 21944 50080 21953
rect 49752 21904 49794 21944
rect 49834 21904 49876 21944
rect 49916 21904 49958 21944
rect 49998 21904 50040 21944
rect 49712 21895 50080 21904
rect 64832 21944 65200 21953
rect 64872 21904 64914 21944
rect 64954 21904 64996 21944
rect 65036 21904 65078 21944
rect 65118 21904 65160 21944
rect 64832 21895 65200 21904
rect 79952 21944 80320 21953
rect 79992 21904 80034 21944
rect 80074 21904 80116 21944
rect 80156 21904 80198 21944
rect 80238 21904 80280 21944
rect 79952 21895 80320 21904
rect 95072 21944 95440 21953
rect 95112 21904 95154 21944
rect 95194 21904 95236 21944
rect 95276 21904 95318 21944
rect 95358 21904 95400 21944
rect 95072 21895 95440 21904
rect 3112 21188 3480 21197
rect 3152 21148 3194 21188
rect 3234 21148 3276 21188
rect 3316 21148 3358 21188
rect 3398 21148 3440 21188
rect 3112 21139 3480 21148
rect 18232 21188 18600 21197
rect 18272 21148 18314 21188
rect 18354 21148 18396 21188
rect 18436 21148 18478 21188
rect 18518 21148 18560 21188
rect 18232 21139 18600 21148
rect 33352 21188 33720 21197
rect 33392 21148 33434 21188
rect 33474 21148 33516 21188
rect 33556 21148 33598 21188
rect 33638 21148 33680 21188
rect 33352 21139 33720 21148
rect 48472 21188 48840 21197
rect 48512 21148 48554 21188
rect 48594 21148 48636 21188
rect 48676 21148 48718 21188
rect 48758 21148 48800 21188
rect 48472 21139 48840 21148
rect 63592 21188 63960 21197
rect 63632 21148 63674 21188
rect 63714 21148 63756 21188
rect 63796 21148 63838 21188
rect 63878 21148 63920 21188
rect 63592 21139 63960 21148
rect 78712 21188 79080 21197
rect 78752 21148 78794 21188
rect 78834 21148 78876 21188
rect 78916 21148 78958 21188
rect 78998 21148 79040 21188
rect 78712 21139 79080 21148
rect 93832 21188 94200 21197
rect 93872 21148 93914 21188
rect 93954 21148 93996 21188
rect 94036 21148 94078 21188
rect 94118 21148 94160 21188
rect 93832 21139 94200 21148
rect 4352 20432 4720 20441
rect 4392 20392 4434 20432
rect 4474 20392 4516 20432
rect 4556 20392 4598 20432
rect 4638 20392 4680 20432
rect 4352 20383 4720 20392
rect 19472 20432 19840 20441
rect 19512 20392 19554 20432
rect 19594 20392 19636 20432
rect 19676 20392 19718 20432
rect 19758 20392 19800 20432
rect 19472 20383 19840 20392
rect 34592 20432 34960 20441
rect 34632 20392 34674 20432
rect 34714 20392 34756 20432
rect 34796 20392 34838 20432
rect 34878 20392 34920 20432
rect 34592 20383 34960 20392
rect 49712 20432 50080 20441
rect 49752 20392 49794 20432
rect 49834 20392 49876 20432
rect 49916 20392 49958 20432
rect 49998 20392 50040 20432
rect 49712 20383 50080 20392
rect 64832 20432 65200 20441
rect 64872 20392 64914 20432
rect 64954 20392 64996 20432
rect 65036 20392 65078 20432
rect 65118 20392 65160 20432
rect 64832 20383 65200 20392
rect 79952 20432 80320 20441
rect 79992 20392 80034 20432
rect 80074 20392 80116 20432
rect 80156 20392 80198 20432
rect 80238 20392 80280 20432
rect 79952 20383 80320 20392
rect 95072 20432 95440 20441
rect 95112 20392 95154 20432
rect 95194 20392 95236 20432
rect 95276 20392 95318 20432
rect 95358 20392 95400 20432
rect 95072 20383 95440 20392
rect 3112 19676 3480 19685
rect 3152 19636 3194 19676
rect 3234 19636 3276 19676
rect 3316 19636 3358 19676
rect 3398 19636 3440 19676
rect 3112 19627 3480 19636
rect 18232 19676 18600 19685
rect 18272 19636 18314 19676
rect 18354 19636 18396 19676
rect 18436 19636 18478 19676
rect 18518 19636 18560 19676
rect 18232 19627 18600 19636
rect 33352 19676 33720 19685
rect 33392 19636 33434 19676
rect 33474 19636 33516 19676
rect 33556 19636 33598 19676
rect 33638 19636 33680 19676
rect 33352 19627 33720 19636
rect 48472 19676 48840 19685
rect 48512 19636 48554 19676
rect 48594 19636 48636 19676
rect 48676 19636 48718 19676
rect 48758 19636 48800 19676
rect 48472 19627 48840 19636
rect 63592 19676 63960 19685
rect 63632 19636 63674 19676
rect 63714 19636 63756 19676
rect 63796 19636 63838 19676
rect 63878 19636 63920 19676
rect 63592 19627 63960 19636
rect 78712 19676 79080 19685
rect 78752 19636 78794 19676
rect 78834 19636 78876 19676
rect 78916 19636 78958 19676
rect 78998 19636 79040 19676
rect 78712 19627 79080 19636
rect 93832 19676 94200 19685
rect 93872 19636 93914 19676
rect 93954 19636 93996 19676
rect 94036 19636 94078 19676
rect 94118 19636 94160 19676
rect 93832 19627 94200 19636
rect 4352 18920 4720 18929
rect 4392 18880 4434 18920
rect 4474 18880 4516 18920
rect 4556 18880 4598 18920
rect 4638 18880 4680 18920
rect 4352 18871 4720 18880
rect 19472 18920 19840 18929
rect 19512 18880 19554 18920
rect 19594 18880 19636 18920
rect 19676 18880 19718 18920
rect 19758 18880 19800 18920
rect 19472 18871 19840 18880
rect 34592 18920 34960 18929
rect 34632 18880 34674 18920
rect 34714 18880 34756 18920
rect 34796 18880 34838 18920
rect 34878 18880 34920 18920
rect 34592 18871 34960 18880
rect 49712 18920 50080 18929
rect 49752 18880 49794 18920
rect 49834 18880 49876 18920
rect 49916 18880 49958 18920
rect 49998 18880 50040 18920
rect 49712 18871 50080 18880
rect 64832 18920 65200 18929
rect 64872 18880 64914 18920
rect 64954 18880 64996 18920
rect 65036 18880 65078 18920
rect 65118 18880 65160 18920
rect 64832 18871 65200 18880
rect 79952 18920 80320 18929
rect 79992 18880 80034 18920
rect 80074 18880 80116 18920
rect 80156 18880 80198 18920
rect 80238 18880 80280 18920
rect 79952 18871 80320 18880
rect 95072 18920 95440 18929
rect 95112 18880 95154 18920
rect 95194 18880 95236 18920
rect 95276 18880 95318 18920
rect 95358 18880 95400 18920
rect 95072 18871 95440 18880
rect 3112 18164 3480 18173
rect 3152 18124 3194 18164
rect 3234 18124 3276 18164
rect 3316 18124 3358 18164
rect 3398 18124 3440 18164
rect 3112 18115 3480 18124
rect 18232 18164 18600 18173
rect 18272 18124 18314 18164
rect 18354 18124 18396 18164
rect 18436 18124 18478 18164
rect 18518 18124 18560 18164
rect 18232 18115 18600 18124
rect 33352 18164 33720 18173
rect 33392 18124 33434 18164
rect 33474 18124 33516 18164
rect 33556 18124 33598 18164
rect 33638 18124 33680 18164
rect 33352 18115 33720 18124
rect 48472 18164 48840 18173
rect 48512 18124 48554 18164
rect 48594 18124 48636 18164
rect 48676 18124 48718 18164
rect 48758 18124 48800 18164
rect 48472 18115 48840 18124
rect 63592 18164 63960 18173
rect 63632 18124 63674 18164
rect 63714 18124 63756 18164
rect 63796 18124 63838 18164
rect 63878 18124 63920 18164
rect 63592 18115 63960 18124
rect 78712 18164 79080 18173
rect 78752 18124 78794 18164
rect 78834 18124 78876 18164
rect 78916 18124 78958 18164
rect 78998 18124 79040 18164
rect 78712 18115 79080 18124
rect 93832 18164 94200 18173
rect 93872 18124 93914 18164
rect 93954 18124 93996 18164
rect 94036 18124 94078 18164
rect 94118 18124 94160 18164
rect 93832 18115 94200 18124
rect 4352 17408 4720 17417
rect 4392 17368 4434 17408
rect 4474 17368 4516 17408
rect 4556 17368 4598 17408
rect 4638 17368 4680 17408
rect 4352 17359 4720 17368
rect 19472 17408 19840 17417
rect 19512 17368 19554 17408
rect 19594 17368 19636 17408
rect 19676 17368 19718 17408
rect 19758 17368 19800 17408
rect 19472 17359 19840 17368
rect 34592 17408 34960 17417
rect 34632 17368 34674 17408
rect 34714 17368 34756 17408
rect 34796 17368 34838 17408
rect 34878 17368 34920 17408
rect 34592 17359 34960 17368
rect 49712 17408 50080 17417
rect 49752 17368 49794 17408
rect 49834 17368 49876 17408
rect 49916 17368 49958 17408
rect 49998 17368 50040 17408
rect 49712 17359 50080 17368
rect 64832 17408 65200 17417
rect 64872 17368 64914 17408
rect 64954 17368 64996 17408
rect 65036 17368 65078 17408
rect 65118 17368 65160 17408
rect 64832 17359 65200 17368
rect 79952 17408 80320 17417
rect 79992 17368 80034 17408
rect 80074 17368 80116 17408
rect 80156 17368 80198 17408
rect 80238 17368 80280 17408
rect 79952 17359 80320 17368
rect 95072 17408 95440 17417
rect 95112 17368 95154 17408
rect 95194 17368 95236 17408
rect 95276 17368 95318 17408
rect 95358 17368 95400 17408
rect 95072 17359 95440 17368
rect 3112 16652 3480 16661
rect 3152 16612 3194 16652
rect 3234 16612 3276 16652
rect 3316 16612 3358 16652
rect 3398 16612 3440 16652
rect 3112 16603 3480 16612
rect 18232 16652 18600 16661
rect 18272 16612 18314 16652
rect 18354 16612 18396 16652
rect 18436 16612 18478 16652
rect 18518 16612 18560 16652
rect 18232 16603 18600 16612
rect 33352 16652 33720 16661
rect 33392 16612 33434 16652
rect 33474 16612 33516 16652
rect 33556 16612 33598 16652
rect 33638 16612 33680 16652
rect 33352 16603 33720 16612
rect 48472 16652 48840 16661
rect 48512 16612 48554 16652
rect 48594 16612 48636 16652
rect 48676 16612 48718 16652
rect 48758 16612 48800 16652
rect 48472 16603 48840 16612
rect 63592 16652 63960 16661
rect 63632 16612 63674 16652
rect 63714 16612 63756 16652
rect 63796 16612 63838 16652
rect 63878 16612 63920 16652
rect 63592 16603 63960 16612
rect 78712 16652 79080 16661
rect 78752 16612 78794 16652
rect 78834 16612 78876 16652
rect 78916 16612 78958 16652
rect 78998 16612 79040 16652
rect 78712 16603 79080 16612
rect 93832 16652 94200 16661
rect 93872 16612 93914 16652
rect 93954 16612 93996 16652
rect 94036 16612 94078 16652
rect 94118 16612 94160 16652
rect 93832 16603 94200 16612
rect 4352 15896 4720 15905
rect 4392 15856 4434 15896
rect 4474 15856 4516 15896
rect 4556 15856 4598 15896
rect 4638 15856 4680 15896
rect 4352 15847 4720 15856
rect 19472 15896 19840 15905
rect 19512 15856 19554 15896
rect 19594 15856 19636 15896
rect 19676 15856 19718 15896
rect 19758 15856 19800 15896
rect 19472 15847 19840 15856
rect 34592 15896 34960 15905
rect 34632 15856 34674 15896
rect 34714 15856 34756 15896
rect 34796 15856 34838 15896
rect 34878 15856 34920 15896
rect 34592 15847 34960 15856
rect 49712 15896 50080 15905
rect 49752 15856 49794 15896
rect 49834 15856 49876 15896
rect 49916 15856 49958 15896
rect 49998 15856 50040 15896
rect 49712 15847 50080 15856
rect 64832 15896 65200 15905
rect 64872 15856 64914 15896
rect 64954 15856 64996 15896
rect 65036 15856 65078 15896
rect 65118 15856 65160 15896
rect 64832 15847 65200 15856
rect 79952 15896 80320 15905
rect 79992 15856 80034 15896
rect 80074 15856 80116 15896
rect 80156 15856 80198 15896
rect 80238 15856 80280 15896
rect 79952 15847 80320 15856
rect 95072 15896 95440 15905
rect 95112 15856 95154 15896
rect 95194 15856 95236 15896
rect 95276 15856 95318 15896
rect 95358 15856 95400 15896
rect 95072 15847 95440 15856
rect 3112 15140 3480 15149
rect 3152 15100 3194 15140
rect 3234 15100 3276 15140
rect 3316 15100 3358 15140
rect 3398 15100 3440 15140
rect 3112 15091 3480 15100
rect 18232 15140 18600 15149
rect 18272 15100 18314 15140
rect 18354 15100 18396 15140
rect 18436 15100 18478 15140
rect 18518 15100 18560 15140
rect 18232 15091 18600 15100
rect 33352 15140 33720 15149
rect 33392 15100 33434 15140
rect 33474 15100 33516 15140
rect 33556 15100 33598 15140
rect 33638 15100 33680 15140
rect 33352 15091 33720 15100
rect 48472 15140 48840 15149
rect 48512 15100 48554 15140
rect 48594 15100 48636 15140
rect 48676 15100 48718 15140
rect 48758 15100 48800 15140
rect 48472 15091 48840 15100
rect 63592 15140 63960 15149
rect 63632 15100 63674 15140
rect 63714 15100 63756 15140
rect 63796 15100 63838 15140
rect 63878 15100 63920 15140
rect 63592 15091 63960 15100
rect 78712 15140 79080 15149
rect 78752 15100 78794 15140
rect 78834 15100 78876 15140
rect 78916 15100 78958 15140
rect 78998 15100 79040 15140
rect 78712 15091 79080 15100
rect 93832 15140 94200 15149
rect 93872 15100 93914 15140
rect 93954 15100 93996 15140
rect 94036 15100 94078 15140
rect 94118 15100 94160 15140
rect 93832 15091 94200 15100
rect 4352 14384 4720 14393
rect 4392 14344 4434 14384
rect 4474 14344 4516 14384
rect 4556 14344 4598 14384
rect 4638 14344 4680 14384
rect 4352 14335 4720 14344
rect 19472 14384 19840 14393
rect 19512 14344 19554 14384
rect 19594 14344 19636 14384
rect 19676 14344 19718 14384
rect 19758 14344 19800 14384
rect 19472 14335 19840 14344
rect 34592 14384 34960 14393
rect 34632 14344 34674 14384
rect 34714 14344 34756 14384
rect 34796 14344 34838 14384
rect 34878 14344 34920 14384
rect 34592 14335 34960 14344
rect 49712 14384 50080 14393
rect 49752 14344 49794 14384
rect 49834 14344 49876 14384
rect 49916 14344 49958 14384
rect 49998 14344 50040 14384
rect 49712 14335 50080 14344
rect 64832 14384 65200 14393
rect 64872 14344 64914 14384
rect 64954 14344 64996 14384
rect 65036 14344 65078 14384
rect 65118 14344 65160 14384
rect 64832 14335 65200 14344
rect 79952 14384 80320 14393
rect 79992 14344 80034 14384
rect 80074 14344 80116 14384
rect 80156 14344 80198 14384
rect 80238 14344 80280 14384
rect 79952 14335 80320 14344
rect 95072 14384 95440 14393
rect 95112 14344 95154 14384
rect 95194 14344 95236 14384
rect 95276 14344 95318 14384
rect 95358 14344 95400 14384
rect 95072 14335 95440 14344
rect 3112 13628 3480 13637
rect 3152 13588 3194 13628
rect 3234 13588 3276 13628
rect 3316 13588 3358 13628
rect 3398 13588 3440 13628
rect 3112 13579 3480 13588
rect 18232 13628 18600 13637
rect 18272 13588 18314 13628
rect 18354 13588 18396 13628
rect 18436 13588 18478 13628
rect 18518 13588 18560 13628
rect 18232 13579 18600 13588
rect 33352 13628 33720 13637
rect 33392 13588 33434 13628
rect 33474 13588 33516 13628
rect 33556 13588 33598 13628
rect 33638 13588 33680 13628
rect 33352 13579 33720 13588
rect 48472 13628 48840 13637
rect 48512 13588 48554 13628
rect 48594 13588 48636 13628
rect 48676 13588 48718 13628
rect 48758 13588 48800 13628
rect 48472 13579 48840 13588
rect 63592 13628 63960 13637
rect 63632 13588 63674 13628
rect 63714 13588 63756 13628
rect 63796 13588 63838 13628
rect 63878 13588 63920 13628
rect 63592 13579 63960 13588
rect 78712 13628 79080 13637
rect 78752 13588 78794 13628
rect 78834 13588 78876 13628
rect 78916 13588 78958 13628
rect 78998 13588 79040 13628
rect 78712 13579 79080 13588
rect 93832 13628 94200 13637
rect 93872 13588 93914 13628
rect 93954 13588 93996 13628
rect 94036 13588 94078 13628
rect 94118 13588 94160 13628
rect 93832 13579 94200 13588
rect 4352 12872 4720 12881
rect 4392 12832 4434 12872
rect 4474 12832 4516 12872
rect 4556 12832 4598 12872
rect 4638 12832 4680 12872
rect 4352 12823 4720 12832
rect 19472 12872 19840 12881
rect 19512 12832 19554 12872
rect 19594 12832 19636 12872
rect 19676 12832 19718 12872
rect 19758 12832 19800 12872
rect 19472 12823 19840 12832
rect 34592 12872 34960 12881
rect 34632 12832 34674 12872
rect 34714 12832 34756 12872
rect 34796 12832 34838 12872
rect 34878 12832 34920 12872
rect 34592 12823 34960 12832
rect 49712 12872 50080 12881
rect 49752 12832 49794 12872
rect 49834 12832 49876 12872
rect 49916 12832 49958 12872
rect 49998 12832 50040 12872
rect 49712 12823 50080 12832
rect 64832 12872 65200 12881
rect 64872 12832 64914 12872
rect 64954 12832 64996 12872
rect 65036 12832 65078 12872
rect 65118 12832 65160 12872
rect 64832 12823 65200 12832
rect 79952 12872 80320 12881
rect 79992 12832 80034 12872
rect 80074 12832 80116 12872
rect 80156 12832 80198 12872
rect 80238 12832 80280 12872
rect 79952 12823 80320 12832
rect 95072 12872 95440 12881
rect 95112 12832 95154 12872
rect 95194 12832 95236 12872
rect 95276 12832 95318 12872
rect 95358 12832 95400 12872
rect 95072 12823 95440 12832
rect 3112 12116 3480 12125
rect 3152 12076 3194 12116
rect 3234 12076 3276 12116
rect 3316 12076 3358 12116
rect 3398 12076 3440 12116
rect 3112 12067 3480 12076
rect 18232 12116 18600 12125
rect 18272 12076 18314 12116
rect 18354 12076 18396 12116
rect 18436 12076 18478 12116
rect 18518 12076 18560 12116
rect 18232 12067 18600 12076
rect 33352 12116 33720 12125
rect 33392 12076 33434 12116
rect 33474 12076 33516 12116
rect 33556 12076 33598 12116
rect 33638 12076 33680 12116
rect 33352 12067 33720 12076
rect 48472 12116 48840 12125
rect 48512 12076 48554 12116
rect 48594 12076 48636 12116
rect 48676 12076 48718 12116
rect 48758 12076 48800 12116
rect 48472 12067 48840 12076
rect 63592 12116 63960 12125
rect 63632 12076 63674 12116
rect 63714 12076 63756 12116
rect 63796 12076 63838 12116
rect 63878 12076 63920 12116
rect 63592 12067 63960 12076
rect 78712 12116 79080 12125
rect 78752 12076 78794 12116
rect 78834 12076 78876 12116
rect 78916 12076 78958 12116
rect 78998 12076 79040 12116
rect 78712 12067 79080 12076
rect 93832 12116 94200 12125
rect 93872 12076 93914 12116
rect 93954 12076 93996 12116
rect 94036 12076 94078 12116
rect 94118 12076 94160 12116
rect 93832 12067 94200 12076
rect 4352 11360 4720 11369
rect 4392 11320 4434 11360
rect 4474 11320 4516 11360
rect 4556 11320 4598 11360
rect 4638 11320 4680 11360
rect 4352 11311 4720 11320
rect 19472 11360 19840 11369
rect 19512 11320 19554 11360
rect 19594 11320 19636 11360
rect 19676 11320 19718 11360
rect 19758 11320 19800 11360
rect 19472 11311 19840 11320
rect 34592 11360 34960 11369
rect 34632 11320 34674 11360
rect 34714 11320 34756 11360
rect 34796 11320 34838 11360
rect 34878 11320 34920 11360
rect 34592 11311 34960 11320
rect 49712 11360 50080 11369
rect 49752 11320 49794 11360
rect 49834 11320 49876 11360
rect 49916 11320 49958 11360
rect 49998 11320 50040 11360
rect 49712 11311 50080 11320
rect 64832 11360 65200 11369
rect 64872 11320 64914 11360
rect 64954 11320 64996 11360
rect 65036 11320 65078 11360
rect 65118 11320 65160 11360
rect 64832 11311 65200 11320
rect 79952 11360 80320 11369
rect 79992 11320 80034 11360
rect 80074 11320 80116 11360
rect 80156 11320 80198 11360
rect 80238 11320 80280 11360
rect 79952 11311 80320 11320
rect 95072 11360 95440 11369
rect 95112 11320 95154 11360
rect 95194 11320 95236 11360
rect 95276 11320 95318 11360
rect 95358 11320 95400 11360
rect 95072 11311 95440 11320
rect 3112 10604 3480 10613
rect 3152 10564 3194 10604
rect 3234 10564 3276 10604
rect 3316 10564 3358 10604
rect 3398 10564 3440 10604
rect 3112 10555 3480 10564
rect 18232 10604 18600 10613
rect 18272 10564 18314 10604
rect 18354 10564 18396 10604
rect 18436 10564 18478 10604
rect 18518 10564 18560 10604
rect 18232 10555 18600 10564
rect 33352 10604 33720 10613
rect 33392 10564 33434 10604
rect 33474 10564 33516 10604
rect 33556 10564 33598 10604
rect 33638 10564 33680 10604
rect 33352 10555 33720 10564
rect 48472 10604 48840 10613
rect 48512 10564 48554 10604
rect 48594 10564 48636 10604
rect 48676 10564 48718 10604
rect 48758 10564 48800 10604
rect 48472 10555 48840 10564
rect 63592 10604 63960 10613
rect 63632 10564 63674 10604
rect 63714 10564 63756 10604
rect 63796 10564 63838 10604
rect 63878 10564 63920 10604
rect 63592 10555 63960 10564
rect 78712 10604 79080 10613
rect 78752 10564 78794 10604
rect 78834 10564 78876 10604
rect 78916 10564 78958 10604
rect 78998 10564 79040 10604
rect 78712 10555 79080 10564
rect 93832 10604 94200 10613
rect 93872 10564 93914 10604
rect 93954 10564 93996 10604
rect 94036 10564 94078 10604
rect 94118 10564 94160 10604
rect 93832 10555 94200 10564
rect 4352 9848 4720 9857
rect 4392 9808 4434 9848
rect 4474 9808 4516 9848
rect 4556 9808 4598 9848
rect 4638 9808 4680 9848
rect 4352 9799 4720 9808
rect 19472 9848 19840 9857
rect 19512 9808 19554 9848
rect 19594 9808 19636 9848
rect 19676 9808 19718 9848
rect 19758 9808 19800 9848
rect 19472 9799 19840 9808
rect 34592 9848 34960 9857
rect 34632 9808 34674 9848
rect 34714 9808 34756 9848
rect 34796 9808 34838 9848
rect 34878 9808 34920 9848
rect 34592 9799 34960 9808
rect 49712 9848 50080 9857
rect 49752 9808 49794 9848
rect 49834 9808 49876 9848
rect 49916 9808 49958 9848
rect 49998 9808 50040 9848
rect 49712 9799 50080 9808
rect 64832 9848 65200 9857
rect 64872 9808 64914 9848
rect 64954 9808 64996 9848
rect 65036 9808 65078 9848
rect 65118 9808 65160 9848
rect 64832 9799 65200 9808
rect 79952 9848 80320 9857
rect 79992 9808 80034 9848
rect 80074 9808 80116 9848
rect 80156 9808 80198 9848
rect 80238 9808 80280 9848
rect 79952 9799 80320 9808
rect 95072 9848 95440 9857
rect 95112 9808 95154 9848
rect 95194 9808 95236 9848
rect 95276 9808 95318 9848
rect 95358 9808 95400 9848
rect 95072 9799 95440 9808
rect 3112 9092 3480 9101
rect 3152 9052 3194 9092
rect 3234 9052 3276 9092
rect 3316 9052 3358 9092
rect 3398 9052 3440 9092
rect 3112 9043 3480 9052
rect 18232 9092 18600 9101
rect 18272 9052 18314 9092
rect 18354 9052 18396 9092
rect 18436 9052 18478 9092
rect 18518 9052 18560 9092
rect 18232 9043 18600 9052
rect 33352 9092 33720 9101
rect 33392 9052 33434 9092
rect 33474 9052 33516 9092
rect 33556 9052 33598 9092
rect 33638 9052 33680 9092
rect 33352 9043 33720 9052
rect 48472 9092 48840 9101
rect 48512 9052 48554 9092
rect 48594 9052 48636 9092
rect 48676 9052 48718 9092
rect 48758 9052 48800 9092
rect 48472 9043 48840 9052
rect 63592 9092 63960 9101
rect 63632 9052 63674 9092
rect 63714 9052 63756 9092
rect 63796 9052 63838 9092
rect 63878 9052 63920 9092
rect 63592 9043 63960 9052
rect 78712 9092 79080 9101
rect 78752 9052 78794 9092
rect 78834 9052 78876 9092
rect 78916 9052 78958 9092
rect 78998 9052 79040 9092
rect 78712 9043 79080 9052
rect 93832 9092 94200 9101
rect 93872 9052 93914 9092
rect 93954 9052 93996 9092
rect 94036 9052 94078 9092
rect 94118 9052 94160 9092
rect 93832 9043 94200 9052
rect 4352 8336 4720 8345
rect 4392 8296 4434 8336
rect 4474 8296 4516 8336
rect 4556 8296 4598 8336
rect 4638 8296 4680 8336
rect 4352 8287 4720 8296
rect 19472 8336 19840 8345
rect 19512 8296 19554 8336
rect 19594 8296 19636 8336
rect 19676 8296 19718 8336
rect 19758 8296 19800 8336
rect 19472 8287 19840 8296
rect 34592 8336 34960 8345
rect 34632 8296 34674 8336
rect 34714 8296 34756 8336
rect 34796 8296 34838 8336
rect 34878 8296 34920 8336
rect 34592 8287 34960 8296
rect 49712 8336 50080 8345
rect 49752 8296 49794 8336
rect 49834 8296 49876 8336
rect 49916 8296 49958 8336
rect 49998 8296 50040 8336
rect 49712 8287 50080 8296
rect 64832 8336 65200 8345
rect 64872 8296 64914 8336
rect 64954 8296 64996 8336
rect 65036 8296 65078 8336
rect 65118 8296 65160 8336
rect 64832 8287 65200 8296
rect 79952 8336 80320 8345
rect 79992 8296 80034 8336
rect 80074 8296 80116 8336
rect 80156 8296 80198 8336
rect 80238 8296 80280 8336
rect 79952 8287 80320 8296
rect 95072 8336 95440 8345
rect 95112 8296 95154 8336
rect 95194 8296 95236 8336
rect 95276 8296 95318 8336
rect 95358 8296 95400 8336
rect 95072 8287 95440 8296
rect 3112 7580 3480 7589
rect 3152 7540 3194 7580
rect 3234 7540 3276 7580
rect 3316 7540 3358 7580
rect 3398 7540 3440 7580
rect 3112 7531 3480 7540
rect 18232 7580 18600 7589
rect 18272 7540 18314 7580
rect 18354 7540 18396 7580
rect 18436 7540 18478 7580
rect 18518 7540 18560 7580
rect 18232 7531 18600 7540
rect 33352 7580 33720 7589
rect 33392 7540 33434 7580
rect 33474 7540 33516 7580
rect 33556 7540 33598 7580
rect 33638 7540 33680 7580
rect 33352 7531 33720 7540
rect 48472 7580 48840 7589
rect 48512 7540 48554 7580
rect 48594 7540 48636 7580
rect 48676 7540 48718 7580
rect 48758 7540 48800 7580
rect 48472 7531 48840 7540
rect 63592 7580 63960 7589
rect 63632 7540 63674 7580
rect 63714 7540 63756 7580
rect 63796 7540 63838 7580
rect 63878 7540 63920 7580
rect 63592 7531 63960 7540
rect 78712 7580 79080 7589
rect 78752 7540 78794 7580
rect 78834 7540 78876 7580
rect 78916 7540 78958 7580
rect 78998 7540 79040 7580
rect 78712 7531 79080 7540
rect 93832 7580 94200 7589
rect 93872 7540 93914 7580
rect 93954 7540 93996 7580
rect 94036 7540 94078 7580
rect 94118 7540 94160 7580
rect 93832 7531 94200 7540
rect 4352 6824 4720 6833
rect 4392 6784 4434 6824
rect 4474 6784 4516 6824
rect 4556 6784 4598 6824
rect 4638 6784 4680 6824
rect 4352 6775 4720 6784
rect 19472 6824 19840 6833
rect 19512 6784 19554 6824
rect 19594 6784 19636 6824
rect 19676 6784 19718 6824
rect 19758 6784 19800 6824
rect 19472 6775 19840 6784
rect 34592 6824 34960 6833
rect 34632 6784 34674 6824
rect 34714 6784 34756 6824
rect 34796 6784 34838 6824
rect 34878 6784 34920 6824
rect 34592 6775 34960 6784
rect 49712 6824 50080 6833
rect 49752 6784 49794 6824
rect 49834 6784 49876 6824
rect 49916 6784 49958 6824
rect 49998 6784 50040 6824
rect 49712 6775 50080 6784
rect 64832 6824 65200 6833
rect 64872 6784 64914 6824
rect 64954 6784 64996 6824
rect 65036 6784 65078 6824
rect 65118 6784 65160 6824
rect 64832 6775 65200 6784
rect 79952 6824 80320 6833
rect 79992 6784 80034 6824
rect 80074 6784 80116 6824
rect 80156 6784 80198 6824
rect 80238 6784 80280 6824
rect 79952 6775 80320 6784
rect 95072 6824 95440 6833
rect 95112 6784 95154 6824
rect 95194 6784 95236 6824
rect 95276 6784 95318 6824
rect 95358 6784 95400 6824
rect 95072 6775 95440 6784
rect 3112 6068 3480 6077
rect 3152 6028 3194 6068
rect 3234 6028 3276 6068
rect 3316 6028 3358 6068
rect 3398 6028 3440 6068
rect 3112 6019 3480 6028
rect 18232 6068 18600 6077
rect 18272 6028 18314 6068
rect 18354 6028 18396 6068
rect 18436 6028 18478 6068
rect 18518 6028 18560 6068
rect 18232 6019 18600 6028
rect 33352 6068 33720 6077
rect 33392 6028 33434 6068
rect 33474 6028 33516 6068
rect 33556 6028 33598 6068
rect 33638 6028 33680 6068
rect 33352 6019 33720 6028
rect 48472 6068 48840 6077
rect 48512 6028 48554 6068
rect 48594 6028 48636 6068
rect 48676 6028 48718 6068
rect 48758 6028 48800 6068
rect 48472 6019 48840 6028
rect 63592 6068 63960 6077
rect 63632 6028 63674 6068
rect 63714 6028 63756 6068
rect 63796 6028 63838 6068
rect 63878 6028 63920 6068
rect 63592 6019 63960 6028
rect 78712 6068 79080 6077
rect 78752 6028 78794 6068
rect 78834 6028 78876 6068
rect 78916 6028 78958 6068
rect 78998 6028 79040 6068
rect 78712 6019 79080 6028
rect 93832 6068 94200 6077
rect 93872 6028 93914 6068
rect 93954 6028 93996 6068
rect 94036 6028 94078 6068
rect 94118 6028 94160 6068
rect 93832 6019 94200 6028
rect 4352 5312 4720 5321
rect 4392 5272 4434 5312
rect 4474 5272 4516 5312
rect 4556 5272 4598 5312
rect 4638 5272 4680 5312
rect 4352 5263 4720 5272
rect 19472 5312 19840 5321
rect 19512 5272 19554 5312
rect 19594 5272 19636 5312
rect 19676 5272 19718 5312
rect 19758 5272 19800 5312
rect 19472 5263 19840 5272
rect 34592 5312 34960 5321
rect 34632 5272 34674 5312
rect 34714 5272 34756 5312
rect 34796 5272 34838 5312
rect 34878 5272 34920 5312
rect 34592 5263 34960 5272
rect 49712 5312 50080 5321
rect 49752 5272 49794 5312
rect 49834 5272 49876 5312
rect 49916 5272 49958 5312
rect 49998 5272 50040 5312
rect 49712 5263 50080 5272
rect 64832 5312 65200 5321
rect 64872 5272 64914 5312
rect 64954 5272 64996 5312
rect 65036 5272 65078 5312
rect 65118 5272 65160 5312
rect 64832 5263 65200 5272
rect 79952 5312 80320 5321
rect 79992 5272 80034 5312
rect 80074 5272 80116 5312
rect 80156 5272 80198 5312
rect 80238 5272 80280 5312
rect 79952 5263 80320 5272
rect 95072 5312 95440 5321
rect 95112 5272 95154 5312
rect 95194 5272 95236 5312
rect 95276 5272 95318 5312
rect 95358 5272 95400 5312
rect 95072 5263 95440 5272
rect 3112 4556 3480 4565
rect 3152 4516 3194 4556
rect 3234 4516 3276 4556
rect 3316 4516 3358 4556
rect 3398 4516 3440 4556
rect 3112 4507 3480 4516
rect 18232 4556 18600 4565
rect 18272 4516 18314 4556
rect 18354 4516 18396 4556
rect 18436 4516 18478 4556
rect 18518 4516 18560 4556
rect 18232 4507 18600 4516
rect 33352 4556 33720 4565
rect 33392 4516 33434 4556
rect 33474 4516 33516 4556
rect 33556 4516 33598 4556
rect 33638 4516 33680 4556
rect 33352 4507 33720 4516
rect 48472 4556 48840 4565
rect 48512 4516 48554 4556
rect 48594 4516 48636 4556
rect 48676 4516 48718 4556
rect 48758 4516 48800 4556
rect 48472 4507 48840 4516
rect 63592 4556 63960 4565
rect 63632 4516 63674 4556
rect 63714 4516 63756 4556
rect 63796 4516 63838 4556
rect 63878 4516 63920 4556
rect 63592 4507 63960 4516
rect 78712 4556 79080 4565
rect 78752 4516 78794 4556
rect 78834 4516 78876 4556
rect 78916 4516 78958 4556
rect 78998 4516 79040 4556
rect 78712 4507 79080 4516
rect 93832 4556 94200 4565
rect 93872 4516 93914 4556
rect 93954 4516 93996 4556
rect 94036 4516 94078 4556
rect 94118 4516 94160 4556
rect 93832 4507 94200 4516
rect 4352 3800 4720 3809
rect 4392 3760 4434 3800
rect 4474 3760 4516 3800
rect 4556 3760 4598 3800
rect 4638 3760 4680 3800
rect 4352 3751 4720 3760
rect 19472 3800 19840 3809
rect 19512 3760 19554 3800
rect 19594 3760 19636 3800
rect 19676 3760 19718 3800
rect 19758 3760 19800 3800
rect 19472 3751 19840 3760
rect 34592 3800 34960 3809
rect 34632 3760 34674 3800
rect 34714 3760 34756 3800
rect 34796 3760 34838 3800
rect 34878 3760 34920 3800
rect 34592 3751 34960 3760
rect 49712 3800 50080 3809
rect 49752 3760 49794 3800
rect 49834 3760 49876 3800
rect 49916 3760 49958 3800
rect 49998 3760 50040 3800
rect 49712 3751 50080 3760
rect 64832 3800 65200 3809
rect 64872 3760 64914 3800
rect 64954 3760 64996 3800
rect 65036 3760 65078 3800
rect 65118 3760 65160 3800
rect 64832 3751 65200 3760
rect 79952 3800 80320 3809
rect 79992 3760 80034 3800
rect 80074 3760 80116 3800
rect 80156 3760 80198 3800
rect 80238 3760 80280 3800
rect 79952 3751 80320 3760
rect 95072 3800 95440 3809
rect 95112 3760 95154 3800
rect 95194 3760 95236 3800
rect 95276 3760 95318 3800
rect 95358 3760 95400 3800
rect 95072 3751 95440 3760
rect 3112 3044 3480 3053
rect 3152 3004 3194 3044
rect 3234 3004 3276 3044
rect 3316 3004 3358 3044
rect 3398 3004 3440 3044
rect 3112 2995 3480 3004
rect 18232 3044 18600 3053
rect 18272 3004 18314 3044
rect 18354 3004 18396 3044
rect 18436 3004 18478 3044
rect 18518 3004 18560 3044
rect 18232 2995 18600 3004
rect 33352 3044 33720 3053
rect 33392 3004 33434 3044
rect 33474 3004 33516 3044
rect 33556 3004 33598 3044
rect 33638 3004 33680 3044
rect 33352 2995 33720 3004
rect 48472 3044 48840 3053
rect 48512 3004 48554 3044
rect 48594 3004 48636 3044
rect 48676 3004 48718 3044
rect 48758 3004 48800 3044
rect 48472 2995 48840 3004
rect 63592 3044 63960 3053
rect 63632 3004 63674 3044
rect 63714 3004 63756 3044
rect 63796 3004 63838 3044
rect 63878 3004 63920 3044
rect 63592 2995 63960 3004
rect 78712 3044 79080 3053
rect 78752 3004 78794 3044
rect 78834 3004 78876 3044
rect 78916 3004 78958 3044
rect 78998 3004 79040 3044
rect 78712 2995 79080 3004
rect 93832 3044 94200 3053
rect 93872 3004 93914 3044
rect 93954 3004 93996 3044
rect 94036 3004 94078 3044
rect 94118 3004 94160 3044
rect 93832 2995 94200 3004
rect 4352 2288 4720 2297
rect 4392 2248 4434 2288
rect 4474 2248 4516 2288
rect 4556 2248 4598 2288
rect 4638 2248 4680 2288
rect 4352 2239 4720 2248
rect 19472 2288 19840 2297
rect 19512 2248 19554 2288
rect 19594 2248 19636 2288
rect 19676 2248 19718 2288
rect 19758 2248 19800 2288
rect 19472 2239 19840 2248
rect 34592 2288 34960 2297
rect 34632 2248 34674 2288
rect 34714 2248 34756 2288
rect 34796 2248 34838 2288
rect 34878 2248 34920 2288
rect 34592 2239 34960 2248
rect 49712 2288 50080 2297
rect 49752 2248 49794 2288
rect 49834 2248 49876 2288
rect 49916 2248 49958 2288
rect 49998 2248 50040 2288
rect 49712 2239 50080 2248
rect 64832 2288 65200 2297
rect 64872 2248 64914 2288
rect 64954 2248 64996 2288
rect 65036 2248 65078 2288
rect 65118 2248 65160 2288
rect 64832 2239 65200 2248
rect 79952 2288 80320 2297
rect 79992 2248 80034 2288
rect 80074 2248 80116 2288
rect 80156 2248 80198 2288
rect 80238 2248 80280 2288
rect 79952 2239 80320 2248
rect 95072 2288 95440 2297
rect 95112 2248 95154 2288
rect 95194 2248 95236 2288
rect 95276 2248 95318 2288
rect 95358 2248 95400 2288
rect 95072 2239 95440 2248
rect 3112 1532 3480 1541
rect 3152 1492 3194 1532
rect 3234 1492 3276 1532
rect 3316 1492 3358 1532
rect 3398 1492 3440 1532
rect 3112 1483 3480 1492
rect 18232 1532 18600 1541
rect 18272 1492 18314 1532
rect 18354 1492 18396 1532
rect 18436 1492 18478 1532
rect 18518 1492 18560 1532
rect 18232 1483 18600 1492
rect 33352 1532 33720 1541
rect 33392 1492 33434 1532
rect 33474 1492 33516 1532
rect 33556 1492 33598 1532
rect 33638 1492 33680 1532
rect 33352 1483 33720 1492
rect 48472 1532 48840 1541
rect 48512 1492 48554 1532
rect 48594 1492 48636 1532
rect 48676 1492 48718 1532
rect 48758 1492 48800 1532
rect 48472 1483 48840 1492
rect 63592 1532 63960 1541
rect 63632 1492 63674 1532
rect 63714 1492 63756 1532
rect 63796 1492 63838 1532
rect 63878 1492 63920 1532
rect 63592 1483 63960 1492
rect 78712 1532 79080 1541
rect 78752 1492 78794 1532
rect 78834 1492 78876 1532
rect 78916 1492 78958 1532
rect 78998 1492 79040 1532
rect 78712 1483 79080 1492
rect 93832 1532 94200 1541
rect 93872 1492 93914 1532
rect 93954 1492 93996 1532
rect 94036 1492 94078 1532
rect 94118 1492 94160 1532
rect 93832 1483 94200 1492
rect 4352 776 4720 785
rect 4392 736 4434 776
rect 4474 736 4516 776
rect 4556 736 4598 776
rect 4638 736 4680 776
rect 4352 727 4720 736
rect 19472 776 19840 785
rect 19512 736 19554 776
rect 19594 736 19636 776
rect 19676 736 19718 776
rect 19758 736 19800 776
rect 19472 727 19840 736
rect 34592 776 34960 785
rect 34632 736 34674 776
rect 34714 736 34756 776
rect 34796 736 34838 776
rect 34878 736 34920 776
rect 34592 727 34960 736
rect 49712 776 50080 785
rect 49752 736 49794 776
rect 49834 736 49876 776
rect 49916 736 49958 776
rect 49998 736 50040 776
rect 49712 727 50080 736
rect 64832 776 65200 785
rect 64872 736 64914 776
rect 64954 736 64996 776
rect 65036 736 65078 776
rect 65118 736 65160 776
rect 64832 727 65200 736
rect 79952 776 80320 785
rect 79992 736 80034 776
rect 80074 736 80116 776
rect 80156 736 80198 776
rect 80238 736 80280 776
rect 79952 727 80320 736
rect 95072 776 95440 785
rect 95112 736 95154 776
rect 95194 736 95236 776
rect 95276 736 95318 776
rect 95358 736 95400 776
rect 95072 727 95440 736
<< via4 >>
rect 4352 38536 4392 38576
rect 4434 38536 4474 38576
rect 4516 38536 4556 38576
rect 4598 38536 4638 38576
rect 4680 38536 4720 38576
rect 19472 38536 19512 38576
rect 19554 38536 19594 38576
rect 19636 38536 19676 38576
rect 19718 38536 19758 38576
rect 19800 38536 19840 38576
rect 34592 38536 34632 38576
rect 34674 38536 34714 38576
rect 34756 38536 34796 38576
rect 34838 38536 34878 38576
rect 34920 38536 34960 38576
rect 49712 38536 49752 38576
rect 49794 38536 49834 38576
rect 49876 38536 49916 38576
rect 49958 38536 49998 38576
rect 50040 38536 50080 38576
rect 64832 38536 64872 38576
rect 64914 38536 64954 38576
rect 64996 38536 65036 38576
rect 65078 38536 65118 38576
rect 65160 38536 65200 38576
rect 79952 38536 79992 38576
rect 80034 38536 80074 38576
rect 80116 38536 80156 38576
rect 80198 38536 80238 38576
rect 80280 38536 80320 38576
rect 95072 38536 95112 38576
rect 95154 38536 95194 38576
rect 95236 38536 95276 38576
rect 95318 38536 95358 38576
rect 95400 38536 95440 38576
rect 3112 37780 3152 37820
rect 3194 37780 3234 37820
rect 3276 37780 3316 37820
rect 3358 37780 3398 37820
rect 3440 37780 3480 37820
rect 18232 37780 18272 37820
rect 18314 37780 18354 37820
rect 18396 37780 18436 37820
rect 18478 37780 18518 37820
rect 18560 37780 18600 37820
rect 33352 37780 33392 37820
rect 33434 37780 33474 37820
rect 33516 37780 33556 37820
rect 33598 37780 33638 37820
rect 33680 37780 33720 37820
rect 48472 37780 48512 37820
rect 48554 37780 48594 37820
rect 48636 37780 48676 37820
rect 48718 37780 48758 37820
rect 48800 37780 48840 37820
rect 63592 37780 63632 37820
rect 63674 37780 63714 37820
rect 63756 37780 63796 37820
rect 63838 37780 63878 37820
rect 63920 37780 63960 37820
rect 78712 37780 78752 37820
rect 78794 37780 78834 37820
rect 78876 37780 78916 37820
rect 78958 37780 78998 37820
rect 79040 37780 79080 37820
rect 93832 37780 93872 37820
rect 93914 37780 93954 37820
rect 93996 37780 94036 37820
rect 94078 37780 94118 37820
rect 94160 37780 94200 37820
rect 4352 37024 4392 37064
rect 4434 37024 4474 37064
rect 4516 37024 4556 37064
rect 4598 37024 4638 37064
rect 4680 37024 4720 37064
rect 19472 37024 19512 37064
rect 19554 37024 19594 37064
rect 19636 37024 19676 37064
rect 19718 37024 19758 37064
rect 19800 37024 19840 37064
rect 34592 37024 34632 37064
rect 34674 37024 34714 37064
rect 34756 37024 34796 37064
rect 34838 37024 34878 37064
rect 34920 37024 34960 37064
rect 49712 37024 49752 37064
rect 49794 37024 49834 37064
rect 49876 37024 49916 37064
rect 49958 37024 49998 37064
rect 50040 37024 50080 37064
rect 64832 37024 64872 37064
rect 64914 37024 64954 37064
rect 64996 37024 65036 37064
rect 65078 37024 65118 37064
rect 65160 37024 65200 37064
rect 79952 37024 79992 37064
rect 80034 37024 80074 37064
rect 80116 37024 80156 37064
rect 80198 37024 80238 37064
rect 80280 37024 80320 37064
rect 95072 37024 95112 37064
rect 95154 37024 95194 37064
rect 95236 37024 95276 37064
rect 95318 37024 95358 37064
rect 95400 37024 95440 37064
rect 3112 36268 3152 36308
rect 3194 36268 3234 36308
rect 3276 36268 3316 36308
rect 3358 36268 3398 36308
rect 3440 36268 3480 36308
rect 18232 36268 18272 36308
rect 18314 36268 18354 36308
rect 18396 36268 18436 36308
rect 18478 36268 18518 36308
rect 18560 36268 18600 36308
rect 33352 36268 33392 36308
rect 33434 36268 33474 36308
rect 33516 36268 33556 36308
rect 33598 36268 33638 36308
rect 33680 36268 33720 36308
rect 48472 36268 48512 36308
rect 48554 36268 48594 36308
rect 48636 36268 48676 36308
rect 48718 36268 48758 36308
rect 48800 36268 48840 36308
rect 63592 36268 63632 36308
rect 63674 36268 63714 36308
rect 63756 36268 63796 36308
rect 63838 36268 63878 36308
rect 63920 36268 63960 36308
rect 78712 36268 78752 36308
rect 78794 36268 78834 36308
rect 78876 36268 78916 36308
rect 78958 36268 78998 36308
rect 79040 36268 79080 36308
rect 93832 36268 93872 36308
rect 93914 36268 93954 36308
rect 93996 36268 94036 36308
rect 94078 36268 94118 36308
rect 94160 36268 94200 36308
rect 4352 35512 4392 35552
rect 4434 35512 4474 35552
rect 4516 35512 4556 35552
rect 4598 35512 4638 35552
rect 4680 35512 4720 35552
rect 19472 35512 19512 35552
rect 19554 35512 19594 35552
rect 19636 35512 19676 35552
rect 19718 35512 19758 35552
rect 19800 35512 19840 35552
rect 34592 35512 34632 35552
rect 34674 35512 34714 35552
rect 34756 35512 34796 35552
rect 34838 35512 34878 35552
rect 34920 35512 34960 35552
rect 49712 35512 49752 35552
rect 49794 35512 49834 35552
rect 49876 35512 49916 35552
rect 49958 35512 49998 35552
rect 50040 35512 50080 35552
rect 64832 35512 64872 35552
rect 64914 35512 64954 35552
rect 64996 35512 65036 35552
rect 65078 35512 65118 35552
rect 65160 35512 65200 35552
rect 79952 35512 79992 35552
rect 80034 35512 80074 35552
rect 80116 35512 80156 35552
rect 80198 35512 80238 35552
rect 80280 35512 80320 35552
rect 95072 35512 95112 35552
rect 95154 35512 95194 35552
rect 95236 35512 95276 35552
rect 95318 35512 95358 35552
rect 95400 35512 95440 35552
rect 3112 34756 3152 34796
rect 3194 34756 3234 34796
rect 3276 34756 3316 34796
rect 3358 34756 3398 34796
rect 3440 34756 3480 34796
rect 18232 34756 18272 34796
rect 18314 34756 18354 34796
rect 18396 34756 18436 34796
rect 18478 34756 18518 34796
rect 18560 34756 18600 34796
rect 33352 34756 33392 34796
rect 33434 34756 33474 34796
rect 33516 34756 33556 34796
rect 33598 34756 33638 34796
rect 33680 34756 33720 34796
rect 48472 34756 48512 34796
rect 48554 34756 48594 34796
rect 48636 34756 48676 34796
rect 48718 34756 48758 34796
rect 48800 34756 48840 34796
rect 63592 34756 63632 34796
rect 63674 34756 63714 34796
rect 63756 34756 63796 34796
rect 63838 34756 63878 34796
rect 63920 34756 63960 34796
rect 78712 34756 78752 34796
rect 78794 34756 78834 34796
rect 78876 34756 78916 34796
rect 78958 34756 78998 34796
rect 79040 34756 79080 34796
rect 93832 34756 93872 34796
rect 93914 34756 93954 34796
rect 93996 34756 94036 34796
rect 94078 34756 94118 34796
rect 94160 34756 94200 34796
rect 4352 34000 4392 34040
rect 4434 34000 4474 34040
rect 4516 34000 4556 34040
rect 4598 34000 4638 34040
rect 4680 34000 4720 34040
rect 19472 34000 19512 34040
rect 19554 34000 19594 34040
rect 19636 34000 19676 34040
rect 19718 34000 19758 34040
rect 19800 34000 19840 34040
rect 34592 34000 34632 34040
rect 34674 34000 34714 34040
rect 34756 34000 34796 34040
rect 34838 34000 34878 34040
rect 34920 34000 34960 34040
rect 49712 34000 49752 34040
rect 49794 34000 49834 34040
rect 49876 34000 49916 34040
rect 49958 34000 49998 34040
rect 50040 34000 50080 34040
rect 64832 34000 64872 34040
rect 64914 34000 64954 34040
rect 64996 34000 65036 34040
rect 65078 34000 65118 34040
rect 65160 34000 65200 34040
rect 79952 34000 79992 34040
rect 80034 34000 80074 34040
rect 80116 34000 80156 34040
rect 80198 34000 80238 34040
rect 80280 34000 80320 34040
rect 95072 34000 95112 34040
rect 95154 34000 95194 34040
rect 95236 34000 95276 34040
rect 95318 34000 95358 34040
rect 95400 34000 95440 34040
rect 3112 33244 3152 33284
rect 3194 33244 3234 33284
rect 3276 33244 3316 33284
rect 3358 33244 3398 33284
rect 3440 33244 3480 33284
rect 18232 33244 18272 33284
rect 18314 33244 18354 33284
rect 18396 33244 18436 33284
rect 18478 33244 18518 33284
rect 18560 33244 18600 33284
rect 33352 33244 33392 33284
rect 33434 33244 33474 33284
rect 33516 33244 33556 33284
rect 33598 33244 33638 33284
rect 33680 33244 33720 33284
rect 48472 33244 48512 33284
rect 48554 33244 48594 33284
rect 48636 33244 48676 33284
rect 48718 33244 48758 33284
rect 48800 33244 48840 33284
rect 63592 33244 63632 33284
rect 63674 33244 63714 33284
rect 63756 33244 63796 33284
rect 63838 33244 63878 33284
rect 63920 33244 63960 33284
rect 78712 33244 78752 33284
rect 78794 33244 78834 33284
rect 78876 33244 78916 33284
rect 78958 33244 78998 33284
rect 79040 33244 79080 33284
rect 93832 33244 93872 33284
rect 93914 33244 93954 33284
rect 93996 33244 94036 33284
rect 94078 33244 94118 33284
rect 94160 33244 94200 33284
rect 4352 32488 4392 32528
rect 4434 32488 4474 32528
rect 4516 32488 4556 32528
rect 4598 32488 4638 32528
rect 4680 32488 4720 32528
rect 19472 32488 19512 32528
rect 19554 32488 19594 32528
rect 19636 32488 19676 32528
rect 19718 32488 19758 32528
rect 19800 32488 19840 32528
rect 34592 32488 34632 32528
rect 34674 32488 34714 32528
rect 34756 32488 34796 32528
rect 34838 32488 34878 32528
rect 34920 32488 34960 32528
rect 49712 32488 49752 32528
rect 49794 32488 49834 32528
rect 49876 32488 49916 32528
rect 49958 32488 49998 32528
rect 50040 32488 50080 32528
rect 64832 32488 64872 32528
rect 64914 32488 64954 32528
rect 64996 32488 65036 32528
rect 65078 32488 65118 32528
rect 65160 32488 65200 32528
rect 79952 32488 79992 32528
rect 80034 32488 80074 32528
rect 80116 32488 80156 32528
rect 80198 32488 80238 32528
rect 80280 32488 80320 32528
rect 95072 32488 95112 32528
rect 95154 32488 95194 32528
rect 95236 32488 95276 32528
rect 95318 32488 95358 32528
rect 95400 32488 95440 32528
rect 3112 31732 3152 31772
rect 3194 31732 3234 31772
rect 3276 31732 3316 31772
rect 3358 31732 3398 31772
rect 3440 31732 3480 31772
rect 18232 31732 18272 31772
rect 18314 31732 18354 31772
rect 18396 31732 18436 31772
rect 18478 31732 18518 31772
rect 18560 31732 18600 31772
rect 33352 31732 33392 31772
rect 33434 31732 33474 31772
rect 33516 31732 33556 31772
rect 33598 31732 33638 31772
rect 33680 31732 33720 31772
rect 48472 31732 48512 31772
rect 48554 31732 48594 31772
rect 48636 31732 48676 31772
rect 48718 31732 48758 31772
rect 48800 31732 48840 31772
rect 63592 31732 63632 31772
rect 63674 31732 63714 31772
rect 63756 31732 63796 31772
rect 63838 31732 63878 31772
rect 63920 31732 63960 31772
rect 78712 31732 78752 31772
rect 78794 31732 78834 31772
rect 78876 31732 78916 31772
rect 78958 31732 78998 31772
rect 79040 31732 79080 31772
rect 93832 31732 93872 31772
rect 93914 31732 93954 31772
rect 93996 31732 94036 31772
rect 94078 31732 94118 31772
rect 94160 31732 94200 31772
rect 4352 30976 4392 31016
rect 4434 30976 4474 31016
rect 4516 30976 4556 31016
rect 4598 30976 4638 31016
rect 4680 30976 4720 31016
rect 19472 30976 19512 31016
rect 19554 30976 19594 31016
rect 19636 30976 19676 31016
rect 19718 30976 19758 31016
rect 19800 30976 19840 31016
rect 34592 30976 34632 31016
rect 34674 30976 34714 31016
rect 34756 30976 34796 31016
rect 34838 30976 34878 31016
rect 34920 30976 34960 31016
rect 49712 30976 49752 31016
rect 49794 30976 49834 31016
rect 49876 30976 49916 31016
rect 49958 30976 49998 31016
rect 50040 30976 50080 31016
rect 64832 30976 64872 31016
rect 64914 30976 64954 31016
rect 64996 30976 65036 31016
rect 65078 30976 65118 31016
rect 65160 30976 65200 31016
rect 79952 30976 79992 31016
rect 80034 30976 80074 31016
rect 80116 30976 80156 31016
rect 80198 30976 80238 31016
rect 80280 30976 80320 31016
rect 95072 30976 95112 31016
rect 95154 30976 95194 31016
rect 95236 30976 95276 31016
rect 95318 30976 95358 31016
rect 95400 30976 95440 31016
rect 3112 30220 3152 30260
rect 3194 30220 3234 30260
rect 3276 30220 3316 30260
rect 3358 30220 3398 30260
rect 3440 30220 3480 30260
rect 18232 30220 18272 30260
rect 18314 30220 18354 30260
rect 18396 30220 18436 30260
rect 18478 30220 18518 30260
rect 18560 30220 18600 30260
rect 33352 30220 33392 30260
rect 33434 30220 33474 30260
rect 33516 30220 33556 30260
rect 33598 30220 33638 30260
rect 33680 30220 33720 30260
rect 48472 30220 48512 30260
rect 48554 30220 48594 30260
rect 48636 30220 48676 30260
rect 48718 30220 48758 30260
rect 48800 30220 48840 30260
rect 63592 30220 63632 30260
rect 63674 30220 63714 30260
rect 63756 30220 63796 30260
rect 63838 30220 63878 30260
rect 63920 30220 63960 30260
rect 78712 30220 78752 30260
rect 78794 30220 78834 30260
rect 78876 30220 78916 30260
rect 78958 30220 78998 30260
rect 79040 30220 79080 30260
rect 93832 30220 93872 30260
rect 93914 30220 93954 30260
rect 93996 30220 94036 30260
rect 94078 30220 94118 30260
rect 94160 30220 94200 30260
rect 4352 29464 4392 29504
rect 4434 29464 4474 29504
rect 4516 29464 4556 29504
rect 4598 29464 4638 29504
rect 4680 29464 4720 29504
rect 19472 29464 19512 29504
rect 19554 29464 19594 29504
rect 19636 29464 19676 29504
rect 19718 29464 19758 29504
rect 19800 29464 19840 29504
rect 34592 29464 34632 29504
rect 34674 29464 34714 29504
rect 34756 29464 34796 29504
rect 34838 29464 34878 29504
rect 34920 29464 34960 29504
rect 49712 29464 49752 29504
rect 49794 29464 49834 29504
rect 49876 29464 49916 29504
rect 49958 29464 49998 29504
rect 50040 29464 50080 29504
rect 64832 29464 64872 29504
rect 64914 29464 64954 29504
rect 64996 29464 65036 29504
rect 65078 29464 65118 29504
rect 65160 29464 65200 29504
rect 79952 29464 79992 29504
rect 80034 29464 80074 29504
rect 80116 29464 80156 29504
rect 80198 29464 80238 29504
rect 80280 29464 80320 29504
rect 95072 29464 95112 29504
rect 95154 29464 95194 29504
rect 95236 29464 95276 29504
rect 95318 29464 95358 29504
rect 95400 29464 95440 29504
rect 3112 28708 3152 28748
rect 3194 28708 3234 28748
rect 3276 28708 3316 28748
rect 3358 28708 3398 28748
rect 3440 28708 3480 28748
rect 18232 28708 18272 28748
rect 18314 28708 18354 28748
rect 18396 28708 18436 28748
rect 18478 28708 18518 28748
rect 18560 28708 18600 28748
rect 33352 28708 33392 28748
rect 33434 28708 33474 28748
rect 33516 28708 33556 28748
rect 33598 28708 33638 28748
rect 33680 28708 33720 28748
rect 48472 28708 48512 28748
rect 48554 28708 48594 28748
rect 48636 28708 48676 28748
rect 48718 28708 48758 28748
rect 48800 28708 48840 28748
rect 63592 28708 63632 28748
rect 63674 28708 63714 28748
rect 63756 28708 63796 28748
rect 63838 28708 63878 28748
rect 63920 28708 63960 28748
rect 78712 28708 78752 28748
rect 78794 28708 78834 28748
rect 78876 28708 78916 28748
rect 78958 28708 78998 28748
rect 79040 28708 79080 28748
rect 93832 28708 93872 28748
rect 93914 28708 93954 28748
rect 93996 28708 94036 28748
rect 94078 28708 94118 28748
rect 94160 28708 94200 28748
rect 4352 27952 4392 27992
rect 4434 27952 4474 27992
rect 4516 27952 4556 27992
rect 4598 27952 4638 27992
rect 4680 27952 4720 27992
rect 19472 27952 19512 27992
rect 19554 27952 19594 27992
rect 19636 27952 19676 27992
rect 19718 27952 19758 27992
rect 19800 27952 19840 27992
rect 34592 27952 34632 27992
rect 34674 27952 34714 27992
rect 34756 27952 34796 27992
rect 34838 27952 34878 27992
rect 34920 27952 34960 27992
rect 49712 27952 49752 27992
rect 49794 27952 49834 27992
rect 49876 27952 49916 27992
rect 49958 27952 49998 27992
rect 50040 27952 50080 27992
rect 64832 27952 64872 27992
rect 64914 27952 64954 27992
rect 64996 27952 65036 27992
rect 65078 27952 65118 27992
rect 65160 27952 65200 27992
rect 79952 27952 79992 27992
rect 80034 27952 80074 27992
rect 80116 27952 80156 27992
rect 80198 27952 80238 27992
rect 80280 27952 80320 27992
rect 95072 27952 95112 27992
rect 95154 27952 95194 27992
rect 95236 27952 95276 27992
rect 95318 27952 95358 27992
rect 95400 27952 95440 27992
rect 3112 27196 3152 27236
rect 3194 27196 3234 27236
rect 3276 27196 3316 27236
rect 3358 27196 3398 27236
rect 3440 27196 3480 27236
rect 18232 27196 18272 27236
rect 18314 27196 18354 27236
rect 18396 27196 18436 27236
rect 18478 27196 18518 27236
rect 18560 27196 18600 27236
rect 33352 27196 33392 27236
rect 33434 27196 33474 27236
rect 33516 27196 33556 27236
rect 33598 27196 33638 27236
rect 33680 27196 33720 27236
rect 48472 27196 48512 27236
rect 48554 27196 48594 27236
rect 48636 27196 48676 27236
rect 48718 27196 48758 27236
rect 48800 27196 48840 27236
rect 63592 27196 63632 27236
rect 63674 27196 63714 27236
rect 63756 27196 63796 27236
rect 63838 27196 63878 27236
rect 63920 27196 63960 27236
rect 78712 27196 78752 27236
rect 78794 27196 78834 27236
rect 78876 27196 78916 27236
rect 78958 27196 78998 27236
rect 79040 27196 79080 27236
rect 93832 27196 93872 27236
rect 93914 27196 93954 27236
rect 93996 27196 94036 27236
rect 94078 27196 94118 27236
rect 94160 27196 94200 27236
rect 4352 26440 4392 26480
rect 4434 26440 4474 26480
rect 4516 26440 4556 26480
rect 4598 26440 4638 26480
rect 4680 26440 4720 26480
rect 19472 26440 19512 26480
rect 19554 26440 19594 26480
rect 19636 26440 19676 26480
rect 19718 26440 19758 26480
rect 19800 26440 19840 26480
rect 34592 26440 34632 26480
rect 34674 26440 34714 26480
rect 34756 26440 34796 26480
rect 34838 26440 34878 26480
rect 34920 26440 34960 26480
rect 49712 26440 49752 26480
rect 49794 26440 49834 26480
rect 49876 26440 49916 26480
rect 49958 26440 49998 26480
rect 50040 26440 50080 26480
rect 64832 26440 64872 26480
rect 64914 26440 64954 26480
rect 64996 26440 65036 26480
rect 65078 26440 65118 26480
rect 65160 26440 65200 26480
rect 79952 26440 79992 26480
rect 80034 26440 80074 26480
rect 80116 26440 80156 26480
rect 80198 26440 80238 26480
rect 80280 26440 80320 26480
rect 95072 26440 95112 26480
rect 95154 26440 95194 26480
rect 95236 26440 95276 26480
rect 95318 26440 95358 26480
rect 95400 26440 95440 26480
rect 3112 25684 3152 25724
rect 3194 25684 3234 25724
rect 3276 25684 3316 25724
rect 3358 25684 3398 25724
rect 3440 25684 3480 25724
rect 18232 25684 18272 25724
rect 18314 25684 18354 25724
rect 18396 25684 18436 25724
rect 18478 25684 18518 25724
rect 18560 25684 18600 25724
rect 33352 25684 33392 25724
rect 33434 25684 33474 25724
rect 33516 25684 33556 25724
rect 33598 25684 33638 25724
rect 33680 25684 33720 25724
rect 48472 25684 48512 25724
rect 48554 25684 48594 25724
rect 48636 25684 48676 25724
rect 48718 25684 48758 25724
rect 48800 25684 48840 25724
rect 63592 25684 63632 25724
rect 63674 25684 63714 25724
rect 63756 25684 63796 25724
rect 63838 25684 63878 25724
rect 63920 25684 63960 25724
rect 78712 25684 78752 25724
rect 78794 25684 78834 25724
rect 78876 25684 78916 25724
rect 78958 25684 78998 25724
rect 79040 25684 79080 25724
rect 93832 25684 93872 25724
rect 93914 25684 93954 25724
rect 93996 25684 94036 25724
rect 94078 25684 94118 25724
rect 94160 25684 94200 25724
rect 4352 24928 4392 24968
rect 4434 24928 4474 24968
rect 4516 24928 4556 24968
rect 4598 24928 4638 24968
rect 4680 24928 4720 24968
rect 19472 24928 19512 24968
rect 19554 24928 19594 24968
rect 19636 24928 19676 24968
rect 19718 24928 19758 24968
rect 19800 24928 19840 24968
rect 34592 24928 34632 24968
rect 34674 24928 34714 24968
rect 34756 24928 34796 24968
rect 34838 24928 34878 24968
rect 34920 24928 34960 24968
rect 49712 24928 49752 24968
rect 49794 24928 49834 24968
rect 49876 24928 49916 24968
rect 49958 24928 49998 24968
rect 50040 24928 50080 24968
rect 64832 24928 64872 24968
rect 64914 24928 64954 24968
rect 64996 24928 65036 24968
rect 65078 24928 65118 24968
rect 65160 24928 65200 24968
rect 79952 24928 79992 24968
rect 80034 24928 80074 24968
rect 80116 24928 80156 24968
rect 80198 24928 80238 24968
rect 80280 24928 80320 24968
rect 95072 24928 95112 24968
rect 95154 24928 95194 24968
rect 95236 24928 95276 24968
rect 95318 24928 95358 24968
rect 95400 24928 95440 24968
rect 3112 24172 3152 24212
rect 3194 24172 3234 24212
rect 3276 24172 3316 24212
rect 3358 24172 3398 24212
rect 3440 24172 3480 24212
rect 18232 24172 18272 24212
rect 18314 24172 18354 24212
rect 18396 24172 18436 24212
rect 18478 24172 18518 24212
rect 18560 24172 18600 24212
rect 33352 24172 33392 24212
rect 33434 24172 33474 24212
rect 33516 24172 33556 24212
rect 33598 24172 33638 24212
rect 33680 24172 33720 24212
rect 48472 24172 48512 24212
rect 48554 24172 48594 24212
rect 48636 24172 48676 24212
rect 48718 24172 48758 24212
rect 48800 24172 48840 24212
rect 63592 24172 63632 24212
rect 63674 24172 63714 24212
rect 63756 24172 63796 24212
rect 63838 24172 63878 24212
rect 63920 24172 63960 24212
rect 78712 24172 78752 24212
rect 78794 24172 78834 24212
rect 78876 24172 78916 24212
rect 78958 24172 78998 24212
rect 79040 24172 79080 24212
rect 93832 24172 93872 24212
rect 93914 24172 93954 24212
rect 93996 24172 94036 24212
rect 94078 24172 94118 24212
rect 94160 24172 94200 24212
rect 4352 23416 4392 23456
rect 4434 23416 4474 23456
rect 4516 23416 4556 23456
rect 4598 23416 4638 23456
rect 4680 23416 4720 23456
rect 19472 23416 19512 23456
rect 19554 23416 19594 23456
rect 19636 23416 19676 23456
rect 19718 23416 19758 23456
rect 19800 23416 19840 23456
rect 34592 23416 34632 23456
rect 34674 23416 34714 23456
rect 34756 23416 34796 23456
rect 34838 23416 34878 23456
rect 34920 23416 34960 23456
rect 49712 23416 49752 23456
rect 49794 23416 49834 23456
rect 49876 23416 49916 23456
rect 49958 23416 49998 23456
rect 50040 23416 50080 23456
rect 64832 23416 64872 23456
rect 64914 23416 64954 23456
rect 64996 23416 65036 23456
rect 65078 23416 65118 23456
rect 65160 23416 65200 23456
rect 79952 23416 79992 23456
rect 80034 23416 80074 23456
rect 80116 23416 80156 23456
rect 80198 23416 80238 23456
rect 80280 23416 80320 23456
rect 95072 23416 95112 23456
rect 95154 23416 95194 23456
rect 95236 23416 95276 23456
rect 95318 23416 95358 23456
rect 95400 23416 95440 23456
rect 3112 22660 3152 22700
rect 3194 22660 3234 22700
rect 3276 22660 3316 22700
rect 3358 22660 3398 22700
rect 3440 22660 3480 22700
rect 18232 22660 18272 22700
rect 18314 22660 18354 22700
rect 18396 22660 18436 22700
rect 18478 22660 18518 22700
rect 18560 22660 18600 22700
rect 33352 22660 33392 22700
rect 33434 22660 33474 22700
rect 33516 22660 33556 22700
rect 33598 22660 33638 22700
rect 33680 22660 33720 22700
rect 48472 22660 48512 22700
rect 48554 22660 48594 22700
rect 48636 22660 48676 22700
rect 48718 22660 48758 22700
rect 48800 22660 48840 22700
rect 63592 22660 63632 22700
rect 63674 22660 63714 22700
rect 63756 22660 63796 22700
rect 63838 22660 63878 22700
rect 63920 22660 63960 22700
rect 78712 22660 78752 22700
rect 78794 22660 78834 22700
rect 78876 22660 78916 22700
rect 78958 22660 78998 22700
rect 79040 22660 79080 22700
rect 93832 22660 93872 22700
rect 93914 22660 93954 22700
rect 93996 22660 94036 22700
rect 94078 22660 94118 22700
rect 94160 22660 94200 22700
rect 4352 21904 4392 21944
rect 4434 21904 4474 21944
rect 4516 21904 4556 21944
rect 4598 21904 4638 21944
rect 4680 21904 4720 21944
rect 19472 21904 19512 21944
rect 19554 21904 19594 21944
rect 19636 21904 19676 21944
rect 19718 21904 19758 21944
rect 19800 21904 19840 21944
rect 34592 21904 34632 21944
rect 34674 21904 34714 21944
rect 34756 21904 34796 21944
rect 34838 21904 34878 21944
rect 34920 21904 34960 21944
rect 49712 21904 49752 21944
rect 49794 21904 49834 21944
rect 49876 21904 49916 21944
rect 49958 21904 49998 21944
rect 50040 21904 50080 21944
rect 64832 21904 64872 21944
rect 64914 21904 64954 21944
rect 64996 21904 65036 21944
rect 65078 21904 65118 21944
rect 65160 21904 65200 21944
rect 79952 21904 79992 21944
rect 80034 21904 80074 21944
rect 80116 21904 80156 21944
rect 80198 21904 80238 21944
rect 80280 21904 80320 21944
rect 95072 21904 95112 21944
rect 95154 21904 95194 21944
rect 95236 21904 95276 21944
rect 95318 21904 95358 21944
rect 95400 21904 95440 21944
rect 3112 21148 3152 21188
rect 3194 21148 3234 21188
rect 3276 21148 3316 21188
rect 3358 21148 3398 21188
rect 3440 21148 3480 21188
rect 18232 21148 18272 21188
rect 18314 21148 18354 21188
rect 18396 21148 18436 21188
rect 18478 21148 18518 21188
rect 18560 21148 18600 21188
rect 33352 21148 33392 21188
rect 33434 21148 33474 21188
rect 33516 21148 33556 21188
rect 33598 21148 33638 21188
rect 33680 21148 33720 21188
rect 48472 21148 48512 21188
rect 48554 21148 48594 21188
rect 48636 21148 48676 21188
rect 48718 21148 48758 21188
rect 48800 21148 48840 21188
rect 63592 21148 63632 21188
rect 63674 21148 63714 21188
rect 63756 21148 63796 21188
rect 63838 21148 63878 21188
rect 63920 21148 63960 21188
rect 78712 21148 78752 21188
rect 78794 21148 78834 21188
rect 78876 21148 78916 21188
rect 78958 21148 78998 21188
rect 79040 21148 79080 21188
rect 93832 21148 93872 21188
rect 93914 21148 93954 21188
rect 93996 21148 94036 21188
rect 94078 21148 94118 21188
rect 94160 21148 94200 21188
rect 4352 20392 4392 20432
rect 4434 20392 4474 20432
rect 4516 20392 4556 20432
rect 4598 20392 4638 20432
rect 4680 20392 4720 20432
rect 19472 20392 19512 20432
rect 19554 20392 19594 20432
rect 19636 20392 19676 20432
rect 19718 20392 19758 20432
rect 19800 20392 19840 20432
rect 34592 20392 34632 20432
rect 34674 20392 34714 20432
rect 34756 20392 34796 20432
rect 34838 20392 34878 20432
rect 34920 20392 34960 20432
rect 49712 20392 49752 20432
rect 49794 20392 49834 20432
rect 49876 20392 49916 20432
rect 49958 20392 49998 20432
rect 50040 20392 50080 20432
rect 64832 20392 64872 20432
rect 64914 20392 64954 20432
rect 64996 20392 65036 20432
rect 65078 20392 65118 20432
rect 65160 20392 65200 20432
rect 79952 20392 79992 20432
rect 80034 20392 80074 20432
rect 80116 20392 80156 20432
rect 80198 20392 80238 20432
rect 80280 20392 80320 20432
rect 95072 20392 95112 20432
rect 95154 20392 95194 20432
rect 95236 20392 95276 20432
rect 95318 20392 95358 20432
rect 95400 20392 95440 20432
rect 3112 19636 3152 19676
rect 3194 19636 3234 19676
rect 3276 19636 3316 19676
rect 3358 19636 3398 19676
rect 3440 19636 3480 19676
rect 18232 19636 18272 19676
rect 18314 19636 18354 19676
rect 18396 19636 18436 19676
rect 18478 19636 18518 19676
rect 18560 19636 18600 19676
rect 33352 19636 33392 19676
rect 33434 19636 33474 19676
rect 33516 19636 33556 19676
rect 33598 19636 33638 19676
rect 33680 19636 33720 19676
rect 48472 19636 48512 19676
rect 48554 19636 48594 19676
rect 48636 19636 48676 19676
rect 48718 19636 48758 19676
rect 48800 19636 48840 19676
rect 63592 19636 63632 19676
rect 63674 19636 63714 19676
rect 63756 19636 63796 19676
rect 63838 19636 63878 19676
rect 63920 19636 63960 19676
rect 78712 19636 78752 19676
rect 78794 19636 78834 19676
rect 78876 19636 78916 19676
rect 78958 19636 78998 19676
rect 79040 19636 79080 19676
rect 93832 19636 93872 19676
rect 93914 19636 93954 19676
rect 93996 19636 94036 19676
rect 94078 19636 94118 19676
rect 94160 19636 94200 19676
rect 4352 18880 4392 18920
rect 4434 18880 4474 18920
rect 4516 18880 4556 18920
rect 4598 18880 4638 18920
rect 4680 18880 4720 18920
rect 19472 18880 19512 18920
rect 19554 18880 19594 18920
rect 19636 18880 19676 18920
rect 19718 18880 19758 18920
rect 19800 18880 19840 18920
rect 34592 18880 34632 18920
rect 34674 18880 34714 18920
rect 34756 18880 34796 18920
rect 34838 18880 34878 18920
rect 34920 18880 34960 18920
rect 49712 18880 49752 18920
rect 49794 18880 49834 18920
rect 49876 18880 49916 18920
rect 49958 18880 49998 18920
rect 50040 18880 50080 18920
rect 64832 18880 64872 18920
rect 64914 18880 64954 18920
rect 64996 18880 65036 18920
rect 65078 18880 65118 18920
rect 65160 18880 65200 18920
rect 79952 18880 79992 18920
rect 80034 18880 80074 18920
rect 80116 18880 80156 18920
rect 80198 18880 80238 18920
rect 80280 18880 80320 18920
rect 95072 18880 95112 18920
rect 95154 18880 95194 18920
rect 95236 18880 95276 18920
rect 95318 18880 95358 18920
rect 95400 18880 95440 18920
rect 3112 18124 3152 18164
rect 3194 18124 3234 18164
rect 3276 18124 3316 18164
rect 3358 18124 3398 18164
rect 3440 18124 3480 18164
rect 18232 18124 18272 18164
rect 18314 18124 18354 18164
rect 18396 18124 18436 18164
rect 18478 18124 18518 18164
rect 18560 18124 18600 18164
rect 33352 18124 33392 18164
rect 33434 18124 33474 18164
rect 33516 18124 33556 18164
rect 33598 18124 33638 18164
rect 33680 18124 33720 18164
rect 48472 18124 48512 18164
rect 48554 18124 48594 18164
rect 48636 18124 48676 18164
rect 48718 18124 48758 18164
rect 48800 18124 48840 18164
rect 63592 18124 63632 18164
rect 63674 18124 63714 18164
rect 63756 18124 63796 18164
rect 63838 18124 63878 18164
rect 63920 18124 63960 18164
rect 78712 18124 78752 18164
rect 78794 18124 78834 18164
rect 78876 18124 78916 18164
rect 78958 18124 78998 18164
rect 79040 18124 79080 18164
rect 93832 18124 93872 18164
rect 93914 18124 93954 18164
rect 93996 18124 94036 18164
rect 94078 18124 94118 18164
rect 94160 18124 94200 18164
rect 4352 17368 4392 17408
rect 4434 17368 4474 17408
rect 4516 17368 4556 17408
rect 4598 17368 4638 17408
rect 4680 17368 4720 17408
rect 19472 17368 19512 17408
rect 19554 17368 19594 17408
rect 19636 17368 19676 17408
rect 19718 17368 19758 17408
rect 19800 17368 19840 17408
rect 34592 17368 34632 17408
rect 34674 17368 34714 17408
rect 34756 17368 34796 17408
rect 34838 17368 34878 17408
rect 34920 17368 34960 17408
rect 49712 17368 49752 17408
rect 49794 17368 49834 17408
rect 49876 17368 49916 17408
rect 49958 17368 49998 17408
rect 50040 17368 50080 17408
rect 64832 17368 64872 17408
rect 64914 17368 64954 17408
rect 64996 17368 65036 17408
rect 65078 17368 65118 17408
rect 65160 17368 65200 17408
rect 79952 17368 79992 17408
rect 80034 17368 80074 17408
rect 80116 17368 80156 17408
rect 80198 17368 80238 17408
rect 80280 17368 80320 17408
rect 95072 17368 95112 17408
rect 95154 17368 95194 17408
rect 95236 17368 95276 17408
rect 95318 17368 95358 17408
rect 95400 17368 95440 17408
rect 3112 16612 3152 16652
rect 3194 16612 3234 16652
rect 3276 16612 3316 16652
rect 3358 16612 3398 16652
rect 3440 16612 3480 16652
rect 18232 16612 18272 16652
rect 18314 16612 18354 16652
rect 18396 16612 18436 16652
rect 18478 16612 18518 16652
rect 18560 16612 18600 16652
rect 33352 16612 33392 16652
rect 33434 16612 33474 16652
rect 33516 16612 33556 16652
rect 33598 16612 33638 16652
rect 33680 16612 33720 16652
rect 48472 16612 48512 16652
rect 48554 16612 48594 16652
rect 48636 16612 48676 16652
rect 48718 16612 48758 16652
rect 48800 16612 48840 16652
rect 63592 16612 63632 16652
rect 63674 16612 63714 16652
rect 63756 16612 63796 16652
rect 63838 16612 63878 16652
rect 63920 16612 63960 16652
rect 78712 16612 78752 16652
rect 78794 16612 78834 16652
rect 78876 16612 78916 16652
rect 78958 16612 78998 16652
rect 79040 16612 79080 16652
rect 93832 16612 93872 16652
rect 93914 16612 93954 16652
rect 93996 16612 94036 16652
rect 94078 16612 94118 16652
rect 94160 16612 94200 16652
rect 4352 15856 4392 15896
rect 4434 15856 4474 15896
rect 4516 15856 4556 15896
rect 4598 15856 4638 15896
rect 4680 15856 4720 15896
rect 19472 15856 19512 15896
rect 19554 15856 19594 15896
rect 19636 15856 19676 15896
rect 19718 15856 19758 15896
rect 19800 15856 19840 15896
rect 34592 15856 34632 15896
rect 34674 15856 34714 15896
rect 34756 15856 34796 15896
rect 34838 15856 34878 15896
rect 34920 15856 34960 15896
rect 49712 15856 49752 15896
rect 49794 15856 49834 15896
rect 49876 15856 49916 15896
rect 49958 15856 49998 15896
rect 50040 15856 50080 15896
rect 64832 15856 64872 15896
rect 64914 15856 64954 15896
rect 64996 15856 65036 15896
rect 65078 15856 65118 15896
rect 65160 15856 65200 15896
rect 79952 15856 79992 15896
rect 80034 15856 80074 15896
rect 80116 15856 80156 15896
rect 80198 15856 80238 15896
rect 80280 15856 80320 15896
rect 95072 15856 95112 15896
rect 95154 15856 95194 15896
rect 95236 15856 95276 15896
rect 95318 15856 95358 15896
rect 95400 15856 95440 15896
rect 3112 15100 3152 15140
rect 3194 15100 3234 15140
rect 3276 15100 3316 15140
rect 3358 15100 3398 15140
rect 3440 15100 3480 15140
rect 18232 15100 18272 15140
rect 18314 15100 18354 15140
rect 18396 15100 18436 15140
rect 18478 15100 18518 15140
rect 18560 15100 18600 15140
rect 33352 15100 33392 15140
rect 33434 15100 33474 15140
rect 33516 15100 33556 15140
rect 33598 15100 33638 15140
rect 33680 15100 33720 15140
rect 48472 15100 48512 15140
rect 48554 15100 48594 15140
rect 48636 15100 48676 15140
rect 48718 15100 48758 15140
rect 48800 15100 48840 15140
rect 63592 15100 63632 15140
rect 63674 15100 63714 15140
rect 63756 15100 63796 15140
rect 63838 15100 63878 15140
rect 63920 15100 63960 15140
rect 78712 15100 78752 15140
rect 78794 15100 78834 15140
rect 78876 15100 78916 15140
rect 78958 15100 78998 15140
rect 79040 15100 79080 15140
rect 93832 15100 93872 15140
rect 93914 15100 93954 15140
rect 93996 15100 94036 15140
rect 94078 15100 94118 15140
rect 94160 15100 94200 15140
rect 4352 14344 4392 14384
rect 4434 14344 4474 14384
rect 4516 14344 4556 14384
rect 4598 14344 4638 14384
rect 4680 14344 4720 14384
rect 19472 14344 19512 14384
rect 19554 14344 19594 14384
rect 19636 14344 19676 14384
rect 19718 14344 19758 14384
rect 19800 14344 19840 14384
rect 34592 14344 34632 14384
rect 34674 14344 34714 14384
rect 34756 14344 34796 14384
rect 34838 14344 34878 14384
rect 34920 14344 34960 14384
rect 49712 14344 49752 14384
rect 49794 14344 49834 14384
rect 49876 14344 49916 14384
rect 49958 14344 49998 14384
rect 50040 14344 50080 14384
rect 64832 14344 64872 14384
rect 64914 14344 64954 14384
rect 64996 14344 65036 14384
rect 65078 14344 65118 14384
rect 65160 14344 65200 14384
rect 79952 14344 79992 14384
rect 80034 14344 80074 14384
rect 80116 14344 80156 14384
rect 80198 14344 80238 14384
rect 80280 14344 80320 14384
rect 95072 14344 95112 14384
rect 95154 14344 95194 14384
rect 95236 14344 95276 14384
rect 95318 14344 95358 14384
rect 95400 14344 95440 14384
rect 3112 13588 3152 13628
rect 3194 13588 3234 13628
rect 3276 13588 3316 13628
rect 3358 13588 3398 13628
rect 3440 13588 3480 13628
rect 18232 13588 18272 13628
rect 18314 13588 18354 13628
rect 18396 13588 18436 13628
rect 18478 13588 18518 13628
rect 18560 13588 18600 13628
rect 33352 13588 33392 13628
rect 33434 13588 33474 13628
rect 33516 13588 33556 13628
rect 33598 13588 33638 13628
rect 33680 13588 33720 13628
rect 48472 13588 48512 13628
rect 48554 13588 48594 13628
rect 48636 13588 48676 13628
rect 48718 13588 48758 13628
rect 48800 13588 48840 13628
rect 63592 13588 63632 13628
rect 63674 13588 63714 13628
rect 63756 13588 63796 13628
rect 63838 13588 63878 13628
rect 63920 13588 63960 13628
rect 78712 13588 78752 13628
rect 78794 13588 78834 13628
rect 78876 13588 78916 13628
rect 78958 13588 78998 13628
rect 79040 13588 79080 13628
rect 93832 13588 93872 13628
rect 93914 13588 93954 13628
rect 93996 13588 94036 13628
rect 94078 13588 94118 13628
rect 94160 13588 94200 13628
rect 4352 12832 4392 12872
rect 4434 12832 4474 12872
rect 4516 12832 4556 12872
rect 4598 12832 4638 12872
rect 4680 12832 4720 12872
rect 19472 12832 19512 12872
rect 19554 12832 19594 12872
rect 19636 12832 19676 12872
rect 19718 12832 19758 12872
rect 19800 12832 19840 12872
rect 34592 12832 34632 12872
rect 34674 12832 34714 12872
rect 34756 12832 34796 12872
rect 34838 12832 34878 12872
rect 34920 12832 34960 12872
rect 49712 12832 49752 12872
rect 49794 12832 49834 12872
rect 49876 12832 49916 12872
rect 49958 12832 49998 12872
rect 50040 12832 50080 12872
rect 64832 12832 64872 12872
rect 64914 12832 64954 12872
rect 64996 12832 65036 12872
rect 65078 12832 65118 12872
rect 65160 12832 65200 12872
rect 79952 12832 79992 12872
rect 80034 12832 80074 12872
rect 80116 12832 80156 12872
rect 80198 12832 80238 12872
rect 80280 12832 80320 12872
rect 95072 12832 95112 12872
rect 95154 12832 95194 12872
rect 95236 12832 95276 12872
rect 95318 12832 95358 12872
rect 95400 12832 95440 12872
rect 3112 12076 3152 12116
rect 3194 12076 3234 12116
rect 3276 12076 3316 12116
rect 3358 12076 3398 12116
rect 3440 12076 3480 12116
rect 18232 12076 18272 12116
rect 18314 12076 18354 12116
rect 18396 12076 18436 12116
rect 18478 12076 18518 12116
rect 18560 12076 18600 12116
rect 33352 12076 33392 12116
rect 33434 12076 33474 12116
rect 33516 12076 33556 12116
rect 33598 12076 33638 12116
rect 33680 12076 33720 12116
rect 48472 12076 48512 12116
rect 48554 12076 48594 12116
rect 48636 12076 48676 12116
rect 48718 12076 48758 12116
rect 48800 12076 48840 12116
rect 63592 12076 63632 12116
rect 63674 12076 63714 12116
rect 63756 12076 63796 12116
rect 63838 12076 63878 12116
rect 63920 12076 63960 12116
rect 78712 12076 78752 12116
rect 78794 12076 78834 12116
rect 78876 12076 78916 12116
rect 78958 12076 78998 12116
rect 79040 12076 79080 12116
rect 93832 12076 93872 12116
rect 93914 12076 93954 12116
rect 93996 12076 94036 12116
rect 94078 12076 94118 12116
rect 94160 12076 94200 12116
rect 4352 11320 4392 11360
rect 4434 11320 4474 11360
rect 4516 11320 4556 11360
rect 4598 11320 4638 11360
rect 4680 11320 4720 11360
rect 19472 11320 19512 11360
rect 19554 11320 19594 11360
rect 19636 11320 19676 11360
rect 19718 11320 19758 11360
rect 19800 11320 19840 11360
rect 34592 11320 34632 11360
rect 34674 11320 34714 11360
rect 34756 11320 34796 11360
rect 34838 11320 34878 11360
rect 34920 11320 34960 11360
rect 49712 11320 49752 11360
rect 49794 11320 49834 11360
rect 49876 11320 49916 11360
rect 49958 11320 49998 11360
rect 50040 11320 50080 11360
rect 64832 11320 64872 11360
rect 64914 11320 64954 11360
rect 64996 11320 65036 11360
rect 65078 11320 65118 11360
rect 65160 11320 65200 11360
rect 79952 11320 79992 11360
rect 80034 11320 80074 11360
rect 80116 11320 80156 11360
rect 80198 11320 80238 11360
rect 80280 11320 80320 11360
rect 95072 11320 95112 11360
rect 95154 11320 95194 11360
rect 95236 11320 95276 11360
rect 95318 11320 95358 11360
rect 95400 11320 95440 11360
rect 3112 10564 3152 10604
rect 3194 10564 3234 10604
rect 3276 10564 3316 10604
rect 3358 10564 3398 10604
rect 3440 10564 3480 10604
rect 18232 10564 18272 10604
rect 18314 10564 18354 10604
rect 18396 10564 18436 10604
rect 18478 10564 18518 10604
rect 18560 10564 18600 10604
rect 33352 10564 33392 10604
rect 33434 10564 33474 10604
rect 33516 10564 33556 10604
rect 33598 10564 33638 10604
rect 33680 10564 33720 10604
rect 48472 10564 48512 10604
rect 48554 10564 48594 10604
rect 48636 10564 48676 10604
rect 48718 10564 48758 10604
rect 48800 10564 48840 10604
rect 63592 10564 63632 10604
rect 63674 10564 63714 10604
rect 63756 10564 63796 10604
rect 63838 10564 63878 10604
rect 63920 10564 63960 10604
rect 78712 10564 78752 10604
rect 78794 10564 78834 10604
rect 78876 10564 78916 10604
rect 78958 10564 78998 10604
rect 79040 10564 79080 10604
rect 93832 10564 93872 10604
rect 93914 10564 93954 10604
rect 93996 10564 94036 10604
rect 94078 10564 94118 10604
rect 94160 10564 94200 10604
rect 4352 9808 4392 9848
rect 4434 9808 4474 9848
rect 4516 9808 4556 9848
rect 4598 9808 4638 9848
rect 4680 9808 4720 9848
rect 19472 9808 19512 9848
rect 19554 9808 19594 9848
rect 19636 9808 19676 9848
rect 19718 9808 19758 9848
rect 19800 9808 19840 9848
rect 34592 9808 34632 9848
rect 34674 9808 34714 9848
rect 34756 9808 34796 9848
rect 34838 9808 34878 9848
rect 34920 9808 34960 9848
rect 49712 9808 49752 9848
rect 49794 9808 49834 9848
rect 49876 9808 49916 9848
rect 49958 9808 49998 9848
rect 50040 9808 50080 9848
rect 64832 9808 64872 9848
rect 64914 9808 64954 9848
rect 64996 9808 65036 9848
rect 65078 9808 65118 9848
rect 65160 9808 65200 9848
rect 79952 9808 79992 9848
rect 80034 9808 80074 9848
rect 80116 9808 80156 9848
rect 80198 9808 80238 9848
rect 80280 9808 80320 9848
rect 95072 9808 95112 9848
rect 95154 9808 95194 9848
rect 95236 9808 95276 9848
rect 95318 9808 95358 9848
rect 95400 9808 95440 9848
rect 3112 9052 3152 9092
rect 3194 9052 3234 9092
rect 3276 9052 3316 9092
rect 3358 9052 3398 9092
rect 3440 9052 3480 9092
rect 18232 9052 18272 9092
rect 18314 9052 18354 9092
rect 18396 9052 18436 9092
rect 18478 9052 18518 9092
rect 18560 9052 18600 9092
rect 33352 9052 33392 9092
rect 33434 9052 33474 9092
rect 33516 9052 33556 9092
rect 33598 9052 33638 9092
rect 33680 9052 33720 9092
rect 48472 9052 48512 9092
rect 48554 9052 48594 9092
rect 48636 9052 48676 9092
rect 48718 9052 48758 9092
rect 48800 9052 48840 9092
rect 63592 9052 63632 9092
rect 63674 9052 63714 9092
rect 63756 9052 63796 9092
rect 63838 9052 63878 9092
rect 63920 9052 63960 9092
rect 78712 9052 78752 9092
rect 78794 9052 78834 9092
rect 78876 9052 78916 9092
rect 78958 9052 78998 9092
rect 79040 9052 79080 9092
rect 93832 9052 93872 9092
rect 93914 9052 93954 9092
rect 93996 9052 94036 9092
rect 94078 9052 94118 9092
rect 94160 9052 94200 9092
rect 4352 8296 4392 8336
rect 4434 8296 4474 8336
rect 4516 8296 4556 8336
rect 4598 8296 4638 8336
rect 4680 8296 4720 8336
rect 19472 8296 19512 8336
rect 19554 8296 19594 8336
rect 19636 8296 19676 8336
rect 19718 8296 19758 8336
rect 19800 8296 19840 8336
rect 34592 8296 34632 8336
rect 34674 8296 34714 8336
rect 34756 8296 34796 8336
rect 34838 8296 34878 8336
rect 34920 8296 34960 8336
rect 49712 8296 49752 8336
rect 49794 8296 49834 8336
rect 49876 8296 49916 8336
rect 49958 8296 49998 8336
rect 50040 8296 50080 8336
rect 64832 8296 64872 8336
rect 64914 8296 64954 8336
rect 64996 8296 65036 8336
rect 65078 8296 65118 8336
rect 65160 8296 65200 8336
rect 79952 8296 79992 8336
rect 80034 8296 80074 8336
rect 80116 8296 80156 8336
rect 80198 8296 80238 8336
rect 80280 8296 80320 8336
rect 95072 8296 95112 8336
rect 95154 8296 95194 8336
rect 95236 8296 95276 8336
rect 95318 8296 95358 8336
rect 95400 8296 95440 8336
rect 3112 7540 3152 7580
rect 3194 7540 3234 7580
rect 3276 7540 3316 7580
rect 3358 7540 3398 7580
rect 3440 7540 3480 7580
rect 18232 7540 18272 7580
rect 18314 7540 18354 7580
rect 18396 7540 18436 7580
rect 18478 7540 18518 7580
rect 18560 7540 18600 7580
rect 33352 7540 33392 7580
rect 33434 7540 33474 7580
rect 33516 7540 33556 7580
rect 33598 7540 33638 7580
rect 33680 7540 33720 7580
rect 48472 7540 48512 7580
rect 48554 7540 48594 7580
rect 48636 7540 48676 7580
rect 48718 7540 48758 7580
rect 48800 7540 48840 7580
rect 63592 7540 63632 7580
rect 63674 7540 63714 7580
rect 63756 7540 63796 7580
rect 63838 7540 63878 7580
rect 63920 7540 63960 7580
rect 78712 7540 78752 7580
rect 78794 7540 78834 7580
rect 78876 7540 78916 7580
rect 78958 7540 78998 7580
rect 79040 7540 79080 7580
rect 93832 7540 93872 7580
rect 93914 7540 93954 7580
rect 93996 7540 94036 7580
rect 94078 7540 94118 7580
rect 94160 7540 94200 7580
rect 4352 6784 4392 6824
rect 4434 6784 4474 6824
rect 4516 6784 4556 6824
rect 4598 6784 4638 6824
rect 4680 6784 4720 6824
rect 19472 6784 19512 6824
rect 19554 6784 19594 6824
rect 19636 6784 19676 6824
rect 19718 6784 19758 6824
rect 19800 6784 19840 6824
rect 34592 6784 34632 6824
rect 34674 6784 34714 6824
rect 34756 6784 34796 6824
rect 34838 6784 34878 6824
rect 34920 6784 34960 6824
rect 49712 6784 49752 6824
rect 49794 6784 49834 6824
rect 49876 6784 49916 6824
rect 49958 6784 49998 6824
rect 50040 6784 50080 6824
rect 64832 6784 64872 6824
rect 64914 6784 64954 6824
rect 64996 6784 65036 6824
rect 65078 6784 65118 6824
rect 65160 6784 65200 6824
rect 79952 6784 79992 6824
rect 80034 6784 80074 6824
rect 80116 6784 80156 6824
rect 80198 6784 80238 6824
rect 80280 6784 80320 6824
rect 95072 6784 95112 6824
rect 95154 6784 95194 6824
rect 95236 6784 95276 6824
rect 95318 6784 95358 6824
rect 95400 6784 95440 6824
rect 3112 6028 3152 6068
rect 3194 6028 3234 6068
rect 3276 6028 3316 6068
rect 3358 6028 3398 6068
rect 3440 6028 3480 6068
rect 18232 6028 18272 6068
rect 18314 6028 18354 6068
rect 18396 6028 18436 6068
rect 18478 6028 18518 6068
rect 18560 6028 18600 6068
rect 33352 6028 33392 6068
rect 33434 6028 33474 6068
rect 33516 6028 33556 6068
rect 33598 6028 33638 6068
rect 33680 6028 33720 6068
rect 48472 6028 48512 6068
rect 48554 6028 48594 6068
rect 48636 6028 48676 6068
rect 48718 6028 48758 6068
rect 48800 6028 48840 6068
rect 63592 6028 63632 6068
rect 63674 6028 63714 6068
rect 63756 6028 63796 6068
rect 63838 6028 63878 6068
rect 63920 6028 63960 6068
rect 78712 6028 78752 6068
rect 78794 6028 78834 6068
rect 78876 6028 78916 6068
rect 78958 6028 78998 6068
rect 79040 6028 79080 6068
rect 93832 6028 93872 6068
rect 93914 6028 93954 6068
rect 93996 6028 94036 6068
rect 94078 6028 94118 6068
rect 94160 6028 94200 6068
rect 4352 5272 4392 5312
rect 4434 5272 4474 5312
rect 4516 5272 4556 5312
rect 4598 5272 4638 5312
rect 4680 5272 4720 5312
rect 19472 5272 19512 5312
rect 19554 5272 19594 5312
rect 19636 5272 19676 5312
rect 19718 5272 19758 5312
rect 19800 5272 19840 5312
rect 34592 5272 34632 5312
rect 34674 5272 34714 5312
rect 34756 5272 34796 5312
rect 34838 5272 34878 5312
rect 34920 5272 34960 5312
rect 49712 5272 49752 5312
rect 49794 5272 49834 5312
rect 49876 5272 49916 5312
rect 49958 5272 49998 5312
rect 50040 5272 50080 5312
rect 64832 5272 64872 5312
rect 64914 5272 64954 5312
rect 64996 5272 65036 5312
rect 65078 5272 65118 5312
rect 65160 5272 65200 5312
rect 79952 5272 79992 5312
rect 80034 5272 80074 5312
rect 80116 5272 80156 5312
rect 80198 5272 80238 5312
rect 80280 5272 80320 5312
rect 95072 5272 95112 5312
rect 95154 5272 95194 5312
rect 95236 5272 95276 5312
rect 95318 5272 95358 5312
rect 95400 5272 95440 5312
rect 3112 4516 3152 4556
rect 3194 4516 3234 4556
rect 3276 4516 3316 4556
rect 3358 4516 3398 4556
rect 3440 4516 3480 4556
rect 18232 4516 18272 4556
rect 18314 4516 18354 4556
rect 18396 4516 18436 4556
rect 18478 4516 18518 4556
rect 18560 4516 18600 4556
rect 33352 4516 33392 4556
rect 33434 4516 33474 4556
rect 33516 4516 33556 4556
rect 33598 4516 33638 4556
rect 33680 4516 33720 4556
rect 48472 4516 48512 4556
rect 48554 4516 48594 4556
rect 48636 4516 48676 4556
rect 48718 4516 48758 4556
rect 48800 4516 48840 4556
rect 63592 4516 63632 4556
rect 63674 4516 63714 4556
rect 63756 4516 63796 4556
rect 63838 4516 63878 4556
rect 63920 4516 63960 4556
rect 78712 4516 78752 4556
rect 78794 4516 78834 4556
rect 78876 4516 78916 4556
rect 78958 4516 78998 4556
rect 79040 4516 79080 4556
rect 93832 4516 93872 4556
rect 93914 4516 93954 4556
rect 93996 4516 94036 4556
rect 94078 4516 94118 4556
rect 94160 4516 94200 4556
rect 4352 3760 4392 3800
rect 4434 3760 4474 3800
rect 4516 3760 4556 3800
rect 4598 3760 4638 3800
rect 4680 3760 4720 3800
rect 19472 3760 19512 3800
rect 19554 3760 19594 3800
rect 19636 3760 19676 3800
rect 19718 3760 19758 3800
rect 19800 3760 19840 3800
rect 34592 3760 34632 3800
rect 34674 3760 34714 3800
rect 34756 3760 34796 3800
rect 34838 3760 34878 3800
rect 34920 3760 34960 3800
rect 49712 3760 49752 3800
rect 49794 3760 49834 3800
rect 49876 3760 49916 3800
rect 49958 3760 49998 3800
rect 50040 3760 50080 3800
rect 64832 3760 64872 3800
rect 64914 3760 64954 3800
rect 64996 3760 65036 3800
rect 65078 3760 65118 3800
rect 65160 3760 65200 3800
rect 79952 3760 79992 3800
rect 80034 3760 80074 3800
rect 80116 3760 80156 3800
rect 80198 3760 80238 3800
rect 80280 3760 80320 3800
rect 95072 3760 95112 3800
rect 95154 3760 95194 3800
rect 95236 3760 95276 3800
rect 95318 3760 95358 3800
rect 95400 3760 95440 3800
rect 3112 3004 3152 3044
rect 3194 3004 3234 3044
rect 3276 3004 3316 3044
rect 3358 3004 3398 3044
rect 3440 3004 3480 3044
rect 18232 3004 18272 3044
rect 18314 3004 18354 3044
rect 18396 3004 18436 3044
rect 18478 3004 18518 3044
rect 18560 3004 18600 3044
rect 33352 3004 33392 3044
rect 33434 3004 33474 3044
rect 33516 3004 33556 3044
rect 33598 3004 33638 3044
rect 33680 3004 33720 3044
rect 48472 3004 48512 3044
rect 48554 3004 48594 3044
rect 48636 3004 48676 3044
rect 48718 3004 48758 3044
rect 48800 3004 48840 3044
rect 63592 3004 63632 3044
rect 63674 3004 63714 3044
rect 63756 3004 63796 3044
rect 63838 3004 63878 3044
rect 63920 3004 63960 3044
rect 78712 3004 78752 3044
rect 78794 3004 78834 3044
rect 78876 3004 78916 3044
rect 78958 3004 78998 3044
rect 79040 3004 79080 3044
rect 93832 3004 93872 3044
rect 93914 3004 93954 3044
rect 93996 3004 94036 3044
rect 94078 3004 94118 3044
rect 94160 3004 94200 3044
rect 4352 2248 4392 2288
rect 4434 2248 4474 2288
rect 4516 2248 4556 2288
rect 4598 2248 4638 2288
rect 4680 2248 4720 2288
rect 19472 2248 19512 2288
rect 19554 2248 19594 2288
rect 19636 2248 19676 2288
rect 19718 2248 19758 2288
rect 19800 2248 19840 2288
rect 34592 2248 34632 2288
rect 34674 2248 34714 2288
rect 34756 2248 34796 2288
rect 34838 2248 34878 2288
rect 34920 2248 34960 2288
rect 49712 2248 49752 2288
rect 49794 2248 49834 2288
rect 49876 2248 49916 2288
rect 49958 2248 49998 2288
rect 50040 2248 50080 2288
rect 64832 2248 64872 2288
rect 64914 2248 64954 2288
rect 64996 2248 65036 2288
rect 65078 2248 65118 2288
rect 65160 2248 65200 2288
rect 79952 2248 79992 2288
rect 80034 2248 80074 2288
rect 80116 2248 80156 2288
rect 80198 2248 80238 2288
rect 80280 2248 80320 2288
rect 95072 2248 95112 2288
rect 95154 2248 95194 2288
rect 95236 2248 95276 2288
rect 95318 2248 95358 2288
rect 95400 2248 95440 2288
rect 3112 1492 3152 1532
rect 3194 1492 3234 1532
rect 3276 1492 3316 1532
rect 3358 1492 3398 1532
rect 3440 1492 3480 1532
rect 18232 1492 18272 1532
rect 18314 1492 18354 1532
rect 18396 1492 18436 1532
rect 18478 1492 18518 1532
rect 18560 1492 18600 1532
rect 33352 1492 33392 1532
rect 33434 1492 33474 1532
rect 33516 1492 33556 1532
rect 33598 1492 33638 1532
rect 33680 1492 33720 1532
rect 48472 1492 48512 1532
rect 48554 1492 48594 1532
rect 48636 1492 48676 1532
rect 48718 1492 48758 1532
rect 48800 1492 48840 1532
rect 63592 1492 63632 1532
rect 63674 1492 63714 1532
rect 63756 1492 63796 1532
rect 63838 1492 63878 1532
rect 63920 1492 63960 1532
rect 78712 1492 78752 1532
rect 78794 1492 78834 1532
rect 78876 1492 78916 1532
rect 78958 1492 78998 1532
rect 79040 1492 79080 1532
rect 93832 1492 93872 1532
rect 93914 1492 93954 1532
rect 93996 1492 94036 1532
rect 94078 1492 94118 1532
rect 94160 1492 94200 1532
rect 4352 736 4392 776
rect 4434 736 4474 776
rect 4516 736 4556 776
rect 4598 736 4638 776
rect 4680 736 4720 776
rect 19472 736 19512 776
rect 19554 736 19594 776
rect 19636 736 19676 776
rect 19718 736 19758 776
rect 19800 736 19840 776
rect 34592 736 34632 776
rect 34674 736 34714 776
rect 34756 736 34796 776
rect 34838 736 34878 776
rect 34920 736 34960 776
rect 49712 736 49752 776
rect 49794 736 49834 776
rect 49876 736 49916 776
rect 49958 736 49998 776
rect 50040 736 50080 776
rect 64832 736 64872 776
rect 64914 736 64954 776
rect 64996 736 65036 776
rect 65078 736 65118 776
rect 65160 736 65200 776
rect 79952 736 79992 776
rect 80034 736 80074 776
rect 80116 736 80156 776
rect 80198 736 80238 776
rect 80280 736 80320 776
rect 95072 736 95112 776
rect 95154 736 95194 776
rect 95236 736 95276 776
rect 95318 736 95358 776
rect 95400 736 95440 776
<< metal5 >>
rect 4343 38599 4729 38618
rect 4343 38576 4409 38599
rect 4495 38576 4577 38599
rect 4663 38576 4729 38599
rect 4343 38536 4352 38576
rect 4392 38536 4409 38576
rect 4495 38536 4516 38576
rect 4556 38536 4577 38576
rect 4663 38536 4680 38576
rect 4720 38536 4729 38576
rect 4343 38513 4409 38536
rect 4495 38513 4577 38536
rect 4663 38513 4729 38536
rect 4343 38494 4729 38513
rect 19463 38599 19849 38618
rect 19463 38576 19529 38599
rect 19615 38576 19697 38599
rect 19783 38576 19849 38599
rect 19463 38536 19472 38576
rect 19512 38536 19529 38576
rect 19615 38536 19636 38576
rect 19676 38536 19697 38576
rect 19783 38536 19800 38576
rect 19840 38536 19849 38576
rect 19463 38513 19529 38536
rect 19615 38513 19697 38536
rect 19783 38513 19849 38536
rect 19463 38494 19849 38513
rect 34583 38599 34969 38618
rect 34583 38576 34649 38599
rect 34735 38576 34817 38599
rect 34903 38576 34969 38599
rect 34583 38536 34592 38576
rect 34632 38536 34649 38576
rect 34735 38536 34756 38576
rect 34796 38536 34817 38576
rect 34903 38536 34920 38576
rect 34960 38536 34969 38576
rect 34583 38513 34649 38536
rect 34735 38513 34817 38536
rect 34903 38513 34969 38536
rect 34583 38494 34969 38513
rect 49703 38599 50089 38618
rect 49703 38576 49769 38599
rect 49855 38576 49937 38599
rect 50023 38576 50089 38599
rect 49703 38536 49712 38576
rect 49752 38536 49769 38576
rect 49855 38536 49876 38576
rect 49916 38536 49937 38576
rect 50023 38536 50040 38576
rect 50080 38536 50089 38576
rect 49703 38513 49769 38536
rect 49855 38513 49937 38536
rect 50023 38513 50089 38536
rect 49703 38494 50089 38513
rect 64823 38599 65209 38618
rect 64823 38576 64889 38599
rect 64975 38576 65057 38599
rect 65143 38576 65209 38599
rect 64823 38536 64832 38576
rect 64872 38536 64889 38576
rect 64975 38536 64996 38576
rect 65036 38536 65057 38576
rect 65143 38536 65160 38576
rect 65200 38536 65209 38576
rect 64823 38513 64889 38536
rect 64975 38513 65057 38536
rect 65143 38513 65209 38536
rect 64823 38494 65209 38513
rect 79943 38599 80329 38618
rect 79943 38576 80009 38599
rect 80095 38576 80177 38599
rect 80263 38576 80329 38599
rect 79943 38536 79952 38576
rect 79992 38536 80009 38576
rect 80095 38536 80116 38576
rect 80156 38536 80177 38576
rect 80263 38536 80280 38576
rect 80320 38536 80329 38576
rect 79943 38513 80009 38536
rect 80095 38513 80177 38536
rect 80263 38513 80329 38536
rect 79943 38494 80329 38513
rect 95063 38599 95449 38618
rect 95063 38576 95129 38599
rect 95215 38576 95297 38599
rect 95383 38576 95449 38599
rect 95063 38536 95072 38576
rect 95112 38536 95129 38576
rect 95215 38536 95236 38576
rect 95276 38536 95297 38576
rect 95383 38536 95400 38576
rect 95440 38536 95449 38576
rect 95063 38513 95129 38536
rect 95215 38513 95297 38536
rect 95383 38513 95449 38536
rect 95063 38494 95449 38513
rect 3103 37843 3489 37862
rect 3103 37820 3169 37843
rect 3255 37820 3337 37843
rect 3423 37820 3489 37843
rect 3103 37780 3112 37820
rect 3152 37780 3169 37820
rect 3255 37780 3276 37820
rect 3316 37780 3337 37820
rect 3423 37780 3440 37820
rect 3480 37780 3489 37820
rect 3103 37757 3169 37780
rect 3255 37757 3337 37780
rect 3423 37757 3489 37780
rect 3103 37738 3489 37757
rect 18223 37843 18609 37862
rect 18223 37820 18289 37843
rect 18375 37820 18457 37843
rect 18543 37820 18609 37843
rect 18223 37780 18232 37820
rect 18272 37780 18289 37820
rect 18375 37780 18396 37820
rect 18436 37780 18457 37820
rect 18543 37780 18560 37820
rect 18600 37780 18609 37820
rect 18223 37757 18289 37780
rect 18375 37757 18457 37780
rect 18543 37757 18609 37780
rect 18223 37738 18609 37757
rect 33343 37843 33729 37862
rect 33343 37820 33409 37843
rect 33495 37820 33577 37843
rect 33663 37820 33729 37843
rect 33343 37780 33352 37820
rect 33392 37780 33409 37820
rect 33495 37780 33516 37820
rect 33556 37780 33577 37820
rect 33663 37780 33680 37820
rect 33720 37780 33729 37820
rect 33343 37757 33409 37780
rect 33495 37757 33577 37780
rect 33663 37757 33729 37780
rect 33343 37738 33729 37757
rect 48463 37843 48849 37862
rect 48463 37820 48529 37843
rect 48615 37820 48697 37843
rect 48783 37820 48849 37843
rect 48463 37780 48472 37820
rect 48512 37780 48529 37820
rect 48615 37780 48636 37820
rect 48676 37780 48697 37820
rect 48783 37780 48800 37820
rect 48840 37780 48849 37820
rect 48463 37757 48529 37780
rect 48615 37757 48697 37780
rect 48783 37757 48849 37780
rect 48463 37738 48849 37757
rect 63583 37843 63969 37862
rect 63583 37820 63649 37843
rect 63735 37820 63817 37843
rect 63903 37820 63969 37843
rect 63583 37780 63592 37820
rect 63632 37780 63649 37820
rect 63735 37780 63756 37820
rect 63796 37780 63817 37820
rect 63903 37780 63920 37820
rect 63960 37780 63969 37820
rect 63583 37757 63649 37780
rect 63735 37757 63817 37780
rect 63903 37757 63969 37780
rect 63583 37738 63969 37757
rect 78703 37843 79089 37862
rect 78703 37820 78769 37843
rect 78855 37820 78937 37843
rect 79023 37820 79089 37843
rect 78703 37780 78712 37820
rect 78752 37780 78769 37820
rect 78855 37780 78876 37820
rect 78916 37780 78937 37820
rect 79023 37780 79040 37820
rect 79080 37780 79089 37820
rect 78703 37757 78769 37780
rect 78855 37757 78937 37780
rect 79023 37757 79089 37780
rect 78703 37738 79089 37757
rect 93823 37843 94209 37862
rect 93823 37820 93889 37843
rect 93975 37820 94057 37843
rect 94143 37820 94209 37843
rect 93823 37780 93832 37820
rect 93872 37780 93889 37820
rect 93975 37780 93996 37820
rect 94036 37780 94057 37820
rect 94143 37780 94160 37820
rect 94200 37780 94209 37820
rect 93823 37757 93889 37780
rect 93975 37757 94057 37780
rect 94143 37757 94209 37780
rect 93823 37738 94209 37757
rect 4343 37087 4729 37106
rect 4343 37064 4409 37087
rect 4495 37064 4577 37087
rect 4663 37064 4729 37087
rect 4343 37024 4352 37064
rect 4392 37024 4409 37064
rect 4495 37024 4516 37064
rect 4556 37024 4577 37064
rect 4663 37024 4680 37064
rect 4720 37024 4729 37064
rect 4343 37001 4409 37024
rect 4495 37001 4577 37024
rect 4663 37001 4729 37024
rect 4343 36982 4729 37001
rect 19463 37087 19849 37106
rect 19463 37064 19529 37087
rect 19615 37064 19697 37087
rect 19783 37064 19849 37087
rect 19463 37024 19472 37064
rect 19512 37024 19529 37064
rect 19615 37024 19636 37064
rect 19676 37024 19697 37064
rect 19783 37024 19800 37064
rect 19840 37024 19849 37064
rect 19463 37001 19529 37024
rect 19615 37001 19697 37024
rect 19783 37001 19849 37024
rect 19463 36982 19849 37001
rect 34583 37087 34969 37106
rect 34583 37064 34649 37087
rect 34735 37064 34817 37087
rect 34903 37064 34969 37087
rect 34583 37024 34592 37064
rect 34632 37024 34649 37064
rect 34735 37024 34756 37064
rect 34796 37024 34817 37064
rect 34903 37024 34920 37064
rect 34960 37024 34969 37064
rect 34583 37001 34649 37024
rect 34735 37001 34817 37024
rect 34903 37001 34969 37024
rect 34583 36982 34969 37001
rect 49703 37087 50089 37106
rect 49703 37064 49769 37087
rect 49855 37064 49937 37087
rect 50023 37064 50089 37087
rect 49703 37024 49712 37064
rect 49752 37024 49769 37064
rect 49855 37024 49876 37064
rect 49916 37024 49937 37064
rect 50023 37024 50040 37064
rect 50080 37024 50089 37064
rect 49703 37001 49769 37024
rect 49855 37001 49937 37024
rect 50023 37001 50089 37024
rect 49703 36982 50089 37001
rect 64823 37087 65209 37106
rect 64823 37064 64889 37087
rect 64975 37064 65057 37087
rect 65143 37064 65209 37087
rect 64823 37024 64832 37064
rect 64872 37024 64889 37064
rect 64975 37024 64996 37064
rect 65036 37024 65057 37064
rect 65143 37024 65160 37064
rect 65200 37024 65209 37064
rect 64823 37001 64889 37024
rect 64975 37001 65057 37024
rect 65143 37001 65209 37024
rect 64823 36982 65209 37001
rect 79943 37087 80329 37106
rect 79943 37064 80009 37087
rect 80095 37064 80177 37087
rect 80263 37064 80329 37087
rect 79943 37024 79952 37064
rect 79992 37024 80009 37064
rect 80095 37024 80116 37064
rect 80156 37024 80177 37064
rect 80263 37024 80280 37064
rect 80320 37024 80329 37064
rect 79943 37001 80009 37024
rect 80095 37001 80177 37024
rect 80263 37001 80329 37024
rect 79943 36982 80329 37001
rect 95063 37087 95449 37106
rect 95063 37064 95129 37087
rect 95215 37064 95297 37087
rect 95383 37064 95449 37087
rect 95063 37024 95072 37064
rect 95112 37024 95129 37064
rect 95215 37024 95236 37064
rect 95276 37024 95297 37064
rect 95383 37024 95400 37064
rect 95440 37024 95449 37064
rect 95063 37001 95129 37024
rect 95215 37001 95297 37024
rect 95383 37001 95449 37024
rect 95063 36982 95449 37001
rect 3103 36331 3489 36350
rect 3103 36308 3169 36331
rect 3255 36308 3337 36331
rect 3423 36308 3489 36331
rect 3103 36268 3112 36308
rect 3152 36268 3169 36308
rect 3255 36268 3276 36308
rect 3316 36268 3337 36308
rect 3423 36268 3440 36308
rect 3480 36268 3489 36308
rect 3103 36245 3169 36268
rect 3255 36245 3337 36268
rect 3423 36245 3489 36268
rect 3103 36226 3489 36245
rect 18223 36331 18609 36350
rect 18223 36308 18289 36331
rect 18375 36308 18457 36331
rect 18543 36308 18609 36331
rect 18223 36268 18232 36308
rect 18272 36268 18289 36308
rect 18375 36268 18396 36308
rect 18436 36268 18457 36308
rect 18543 36268 18560 36308
rect 18600 36268 18609 36308
rect 18223 36245 18289 36268
rect 18375 36245 18457 36268
rect 18543 36245 18609 36268
rect 18223 36226 18609 36245
rect 33343 36331 33729 36350
rect 33343 36308 33409 36331
rect 33495 36308 33577 36331
rect 33663 36308 33729 36331
rect 33343 36268 33352 36308
rect 33392 36268 33409 36308
rect 33495 36268 33516 36308
rect 33556 36268 33577 36308
rect 33663 36268 33680 36308
rect 33720 36268 33729 36308
rect 33343 36245 33409 36268
rect 33495 36245 33577 36268
rect 33663 36245 33729 36268
rect 33343 36226 33729 36245
rect 48463 36331 48849 36350
rect 48463 36308 48529 36331
rect 48615 36308 48697 36331
rect 48783 36308 48849 36331
rect 48463 36268 48472 36308
rect 48512 36268 48529 36308
rect 48615 36268 48636 36308
rect 48676 36268 48697 36308
rect 48783 36268 48800 36308
rect 48840 36268 48849 36308
rect 48463 36245 48529 36268
rect 48615 36245 48697 36268
rect 48783 36245 48849 36268
rect 48463 36226 48849 36245
rect 63583 36331 63969 36350
rect 63583 36308 63649 36331
rect 63735 36308 63817 36331
rect 63903 36308 63969 36331
rect 63583 36268 63592 36308
rect 63632 36268 63649 36308
rect 63735 36268 63756 36308
rect 63796 36268 63817 36308
rect 63903 36268 63920 36308
rect 63960 36268 63969 36308
rect 63583 36245 63649 36268
rect 63735 36245 63817 36268
rect 63903 36245 63969 36268
rect 63583 36226 63969 36245
rect 78703 36331 79089 36350
rect 78703 36308 78769 36331
rect 78855 36308 78937 36331
rect 79023 36308 79089 36331
rect 78703 36268 78712 36308
rect 78752 36268 78769 36308
rect 78855 36268 78876 36308
rect 78916 36268 78937 36308
rect 79023 36268 79040 36308
rect 79080 36268 79089 36308
rect 78703 36245 78769 36268
rect 78855 36245 78937 36268
rect 79023 36245 79089 36268
rect 78703 36226 79089 36245
rect 93823 36331 94209 36350
rect 93823 36308 93889 36331
rect 93975 36308 94057 36331
rect 94143 36308 94209 36331
rect 93823 36268 93832 36308
rect 93872 36268 93889 36308
rect 93975 36268 93996 36308
rect 94036 36268 94057 36308
rect 94143 36268 94160 36308
rect 94200 36268 94209 36308
rect 93823 36245 93889 36268
rect 93975 36245 94057 36268
rect 94143 36245 94209 36268
rect 93823 36226 94209 36245
rect 4343 35575 4729 35594
rect 4343 35552 4409 35575
rect 4495 35552 4577 35575
rect 4663 35552 4729 35575
rect 4343 35512 4352 35552
rect 4392 35512 4409 35552
rect 4495 35512 4516 35552
rect 4556 35512 4577 35552
rect 4663 35512 4680 35552
rect 4720 35512 4729 35552
rect 4343 35489 4409 35512
rect 4495 35489 4577 35512
rect 4663 35489 4729 35512
rect 4343 35470 4729 35489
rect 19463 35575 19849 35594
rect 19463 35552 19529 35575
rect 19615 35552 19697 35575
rect 19783 35552 19849 35575
rect 19463 35512 19472 35552
rect 19512 35512 19529 35552
rect 19615 35512 19636 35552
rect 19676 35512 19697 35552
rect 19783 35512 19800 35552
rect 19840 35512 19849 35552
rect 19463 35489 19529 35512
rect 19615 35489 19697 35512
rect 19783 35489 19849 35512
rect 19463 35470 19849 35489
rect 34583 35575 34969 35594
rect 34583 35552 34649 35575
rect 34735 35552 34817 35575
rect 34903 35552 34969 35575
rect 34583 35512 34592 35552
rect 34632 35512 34649 35552
rect 34735 35512 34756 35552
rect 34796 35512 34817 35552
rect 34903 35512 34920 35552
rect 34960 35512 34969 35552
rect 34583 35489 34649 35512
rect 34735 35489 34817 35512
rect 34903 35489 34969 35512
rect 34583 35470 34969 35489
rect 49703 35575 50089 35594
rect 49703 35552 49769 35575
rect 49855 35552 49937 35575
rect 50023 35552 50089 35575
rect 49703 35512 49712 35552
rect 49752 35512 49769 35552
rect 49855 35512 49876 35552
rect 49916 35512 49937 35552
rect 50023 35512 50040 35552
rect 50080 35512 50089 35552
rect 49703 35489 49769 35512
rect 49855 35489 49937 35512
rect 50023 35489 50089 35512
rect 49703 35470 50089 35489
rect 64823 35575 65209 35594
rect 64823 35552 64889 35575
rect 64975 35552 65057 35575
rect 65143 35552 65209 35575
rect 64823 35512 64832 35552
rect 64872 35512 64889 35552
rect 64975 35512 64996 35552
rect 65036 35512 65057 35552
rect 65143 35512 65160 35552
rect 65200 35512 65209 35552
rect 64823 35489 64889 35512
rect 64975 35489 65057 35512
rect 65143 35489 65209 35512
rect 64823 35470 65209 35489
rect 79943 35575 80329 35594
rect 79943 35552 80009 35575
rect 80095 35552 80177 35575
rect 80263 35552 80329 35575
rect 79943 35512 79952 35552
rect 79992 35512 80009 35552
rect 80095 35512 80116 35552
rect 80156 35512 80177 35552
rect 80263 35512 80280 35552
rect 80320 35512 80329 35552
rect 79943 35489 80009 35512
rect 80095 35489 80177 35512
rect 80263 35489 80329 35512
rect 79943 35470 80329 35489
rect 95063 35575 95449 35594
rect 95063 35552 95129 35575
rect 95215 35552 95297 35575
rect 95383 35552 95449 35575
rect 95063 35512 95072 35552
rect 95112 35512 95129 35552
rect 95215 35512 95236 35552
rect 95276 35512 95297 35552
rect 95383 35512 95400 35552
rect 95440 35512 95449 35552
rect 95063 35489 95129 35512
rect 95215 35489 95297 35512
rect 95383 35489 95449 35512
rect 95063 35470 95449 35489
rect 3103 34819 3489 34838
rect 3103 34796 3169 34819
rect 3255 34796 3337 34819
rect 3423 34796 3489 34819
rect 3103 34756 3112 34796
rect 3152 34756 3169 34796
rect 3255 34756 3276 34796
rect 3316 34756 3337 34796
rect 3423 34756 3440 34796
rect 3480 34756 3489 34796
rect 3103 34733 3169 34756
rect 3255 34733 3337 34756
rect 3423 34733 3489 34756
rect 3103 34714 3489 34733
rect 18223 34819 18609 34838
rect 18223 34796 18289 34819
rect 18375 34796 18457 34819
rect 18543 34796 18609 34819
rect 18223 34756 18232 34796
rect 18272 34756 18289 34796
rect 18375 34756 18396 34796
rect 18436 34756 18457 34796
rect 18543 34756 18560 34796
rect 18600 34756 18609 34796
rect 18223 34733 18289 34756
rect 18375 34733 18457 34756
rect 18543 34733 18609 34756
rect 18223 34714 18609 34733
rect 33343 34819 33729 34838
rect 33343 34796 33409 34819
rect 33495 34796 33577 34819
rect 33663 34796 33729 34819
rect 33343 34756 33352 34796
rect 33392 34756 33409 34796
rect 33495 34756 33516 34796
rect 33556 34756 33577 34796
rect 33663 34756 33680 34796
rect 33720 34756 33729 34796
rect 33343 34733 33409 34756
rect 33495 34733 33577 34756
rect 33663 34733 33729 34756
rect 33343 34714 33729 34733
rect 48463 34819 48849 34838
rect 48463 34796 48529 34819
rect 48615 34796 48697 34819
rect 48783 34796 48849 34819
rect 48463 34756 48472 34796
rect 48512 34756 48529 34796
rect 48615 34756 48636 34796
rect 48676 34756 48697 34796
rect 48783 34756 48800 34796
rect 48840 34756 48849 34796
rect 48463 34733 48529 34756
rect 48615 34733 48697 34756
rect 48783 34733 48849 34756
rect 48463 34714 48849 34733
rect 63583 34819 63969 34838
rect 63583 34796 63649 34819
rect 63735 34796 63817 34819
rect 63903 34796 63969 34819
rect 63583 34756 63592 34796
rect 63632 34756 63649 34796
rect 63735 34756 63756 34796
rect 63796 34756 63817 34796
rect 63903 34756 63920 34796
rect 63960 34756 63969 34796
rect 63583 34733 63649 34756
rect 63735 34733 63817 34756
rect 63903 34733 63969 34756
rect 63583 34714 63969 34733
rect 78703 34819 79089 34838
rect 78703 34796 78769 34819
rect 78855 34796 78937 34819
rect 79023 34796 79089 34819
rect 78703 34756 78712 34796
rect 78752 34756 78769 34796
rect 78855 34756 78876 34796
rect 78916 34756 78937 34796
rect 79023 34756 79040 34796
rect 79080 34756 79089 34796
rect 78703 34733 78769 34756
rect 78855 34733 78937 34756
rect 79023 34733 79089 34756
rect 78703 34714 79089 34733
rect 93823 34819 94209 34838
rect 93823 34796 93889 34819
rect 93975 34796 94057 34819
rect 94143 34796 94209 34819
rect 93823 34756 93832 34796
rect 93872 34756 93889 34796
rect 93975 34756 93996 34796
rect 94036 34756 94057 34796
rect 94143 34756 94160 34796
rect 94200 34756 94209 34796
rect 93823 34733 93889 34756
rect 93975 34733 94057 34756
rect 94143 34733 94209 34756
rect 93823 34714 94209 34733
rect 4343 34063 4729 34082
rect 4343 34040 4409 34063
rect 4495 34040 4577 34063
rect 4663 34040 4729 34063
rect 4343 34000 4352 34040
rect 4392 34000 4409 34040
rect 4495 34000 4516 34040
rect 4556 34000 4577 34040
rect 4663 34000 4680 34040
rect 4720 34000 4729 34040
rect 4343 33977 4409 34000
rect 4495 33977 4577 34000
rect 4663 33977 4729 34000
rect 4343 33958 4729 33977
rect 19463 34063 19849 34082
rect 19463 34040 19529 34063
rect 19615 34040 19697 34063
rect 19783 34040 19849 34063
rect 19463 34000 19472 34040
rect 19512 34000 19529 34040
rect 19615 34000 19636 34040
rect 19676 34000 19697 34040
rect 19783 34000 19800 34040
rect 19840 34000 19849 34040
rect 19463 33977 19529 34000
rect 19615 33977 19697 34000
rect 19783 33977 19849 34000
rect 19463 33958 19849 33977
rect 34583 34063 34969 34082
rect 34583 34040 34649 34063
rect 34735 34040 34817 34063
rect 34903 34040 34969 34063
rect 34583 34000 34592 34040
rect 34632 34000 34649 34040
rect 34735 34000 34756 34040
rect 34796 34000 34817 34040
rect 34903 34000 34920 34040
rect 34960 34000 34969 34040
rect 34583 33977 34649 34000
rect 34735 33977 34817 34000
rect 34903 33977 34969 34000
rect 34583 33958 34969 33977
rect 49703 34063 50089 34082
rect 49703 34040 49769 34063
rect 49855 34040 49937 34063
rect 50023 34040 50089 34063
rect 49703 34000 49712 34040
rect 49752 34000 49769 34040
rect 49855 34000 49876 34040
rect 49916 34000 49937 34040
rect 50023 34000 50040 34040
rect 50080 34000 50089 34040
rect 49703 33977 49769 34000
rect 49855 33977 49937 34000
rect 50023 33977 50089 34000
rect 49703 33958 50089 33977
rect 64823 34063 65209 34082
rect 64823 34040 64889 34063
rect 64975 34040 65057 34063
rect 65143 34040 65209 34063
rect 64823 34000 64832 34040
rect 64872 34000 64889 34040
rect 64975 34000 64996 34040
rect 65036 34000 65057 34040
rect 65143 34000 65160 34040
rect 65200 34000 65209 34040
rect 64823 33977 64889 34000
rect 64975 33977 65057 34000
rect 65143 33977 65209 34000
rect 64823 33958 65209 33977
rect 79943 34063 80329 34082
rect 79943 34040 80009 34063
rect 80095 34040 80177 34063
rect 80263 34040 80329 34063
rect 79943 34000 79952 34040
rect 79992 34000 80009 34040
rect 80095 34000 80116 34040
rect 80156 34000 80177 34040
rect 80263 34000 80280 34040
rect 80320 34000 80329 34040
rect 79943 33977 80009 34000
rect 80095 33977 80177 34000
rect 80263 33977 80329 34000
rect 79943 33958 80329 33977
rect 95063 34063 95449 34082
rect 95063 34040 95129 34063
rect 95215 34040 95297 34063
rect 95383 34040 95449 34063
rect 95063 34000 95072 34040
rect 95112 34000 95129 34040
rect 95215 34000 95236 34040
rect 95276 34000 95297 34040
rect 95383 34000 95400 34040
rect 95440 34000 95449 34040
rect 95063 33977 95129 34000
rect 95215 33977 95297 34000
rect 95383 33977 95449 34000
rect 95063 33958 95449 33977
rect 3103 33307 3489 33326
rect 3103 33284 3169 33307
rect 3255 33284 3337 33307
rect 3423 33284 3489 33307
rect 3103 33244 3112 33284
rect 3152 33244 3169 33284
rect 3255 33244 3276 33284
rect 3316 33244 3337 33284
rect 3423 33244 3440 33284
rect 3480 33244 3489 33284
rect 3103 33221 3169 33244
rect 3255 33221 3337 33244
rect 3423 33221 3489 33244
rect 3103 33202 3489 33221
rect 18223 33307 18609 33326
rect 18223 33284 18289 33307
rect 18375 33284 18457 33307
rect 18543 33284 18609 33307
rect 18223 33244 18232 33284
rect 18272 33244 18289 33284
rect 18375 33244 18396 33284
rect 18436 33244 18457 33284
rect 18543 33244 18560 33284
rect 18600 33244 18609 33284
rect 18223 33221 18289 33244
rect 18375 33221 18457 33244
rect 18543 33221 18609 33244
rect 18223 33202 18609 33221
rect 33343 33307 33729 33326
rect 33343 33284 33409 33307
rect 33495 33284 33577 33307
rect 33663 33284 33729 33307
rect 33343 33244 33352 33284
rect 33392 33244 33409 33284
rect 33495 33244 33516 33284
rect 33556 33244 33577 33284
rect 33663 33244 33680 33284
rect 33720 33244 33729 33284
rect 33343 33221 33409 33244
rect 33495 33221 33577 33244
rect 33663 33221 33729 33244
rect 33343 33202 33729 33221
rect 48463 33307 48849 33326
rect 48463 33284 48529 33307
rect 48615 33284 48697 33307
rect 48783 33284 48849 33307
rect 48463 33244 48472 33284
rect 48512 33244 48529 33284
rect 48615 33244 48636 33284
rect 48676 33244 48697 33284
rect 48783 33244 48800 33284
rect 48840 33244 48849 33284
rect 48463 33221 48529 33244
rect 48615 33221 48697 33244
rect 48783 33221 48849 33244
rect 48463 33202 48849 33221
rect 63583 33307 63969 33326
rect 63583 33284 63649 33307
rect 63735 33284 63817 33307
rect 63903 33284 63969 33307
rect 63583 33244 63592 33284
rect 63632 33244 63649 33284
rect 63735 33244 63756 33284
rect 63796 33244 63817 33284
rect 63903 33244 63920 33284
rect 63960 33244 63969 33284
rect 63583 33221 63649 33244
rect 63735 33221 63817 33244
rect 63903 33221 63969 33244
rect 63583 33202 63969 33221
rect 78703 33307 79089 33326
rect 78703 33284 78769 33307
rect 78855 33284 78937 33307
rect 79023 33284 79089 33307
rect 78703 33244 78712 33284
rect 78752 33244 78769 33284
rect 78855 33244 78876 33284
rect 78916 33244 78937 33284
rect 79023 33244 79040 33284
rect 79080 33244 79089 33284
rect 78703 33221 78769 33244
rect 78855 33221 78937 33244
rect 79023 33221 79089 33244
rect 78703 33202 79089 33221
rect 93823 33307 94209 33326
rect 93823 33284 93889 33307
rect 93975 33284 94057 33307
rect 94143 33284 94209 33307
rect 93823 33244 93832 33284
rect 93872 33244 93889 33284
rect 93975 33244 93996 33284
rect 94036 33244 94057 33284
rect 94143 33244 94160 33284
rect 94200 33244 94209 33284
rect 93823 33221 93889 33244
rect 93975 33221 94057 33244
rect 94143 33221 94209 33244
rect 93823 33202 94209 33221
rect 4343 32551 4729 32570
rect 4343 32528 4409 32551
rect 4495 32528 4577 32551
rect 4663 32528 4729 32551
rect 4343 32488 4352 32528
rect 4392 32488 4409 32528
rect 4495 32488 4516 32528
rect 4556 32488 4577 32528
rect 4663 32488 4680 32528
rect 4720 32488 4729 32528
rect 4343 32465 4409 32488
rect 4495 32465 4577 32488
rect 4663 32465 4729 32488
rect 4343 32446 4729 32465
rect 19463 32551 19849 32570
rect 19463 32528 19529 32551
rect 19615 32528 19697 32551
rect 19783 32528 19849 32551
rect 19463 32488 19472 32528
rect 19512 32488 19529 32528
rect 19615 32488 19636 32528
rect 19676 32488 19697 32528
rect 19783 32488 19800 32528
rect 19840 32488 19849 32528
rect 19463 32465 19529 32488
rect 19615 32465 19697 32488
rect 19783 32465 19849 32488
rect 19463 32446 19849 32465
rect 34583 32551 34969 32570
rect 34583 32528 34649 32551
rect 34735 32528 34817 32551
rect 34903 32528 34969 32551
rect 34583 32488 34592 32528
rect 34632 32488 34649 32528
rect 34735 32488 34756 32528
rect 34796 32488 34817 32528
rect 34903 32488 34920 32528
rect 34960 32488 34969 32528
rect 34583 32465 34649 32488
rect 34735 32465 34817 32488
rect 34903 32465 34969 32488
rect 34583 32446 34969 32465
rect 49703 32551 50089 32570
rect 49703 32528 49769 32551
rect 49855 32528 49937 32551
rect 50023 32528 50089 32551
rect 49703 32488 49712 32528
rect 49752 32488 49769 32528
rect 49855 32488 49876 32528
rect 49916 32488 49937 32528
rect 50023 32488 50040 32528
rect 50080 32488 50089 32528
rect 49703 32465 49769 32488
rect 49855 32465 49937 32488
rect 50023 32465 50089 32488
rect 49703 32446 50089 32465
rect 64823 32551 65209 32570
rect 64823 32528 64889 32551
rect 64975 32528 65057 32551
rect 65143 32528 65209 32551
rect 64823 32488 64832 32528
rect 64872 32488 64889 32528
rect 64975 32488 64996 32528
rect 65036 32488 65057 32528
rect 65143 32488 65160 32528
rect 65200 32488 65209 32528
rect 64823 32465 64889 32488
rect 64975 32465 65057 32488
rect 65143 32465 65209 32488
rect 64823 32446 65209 32465
rect 79943 32551 80329 32570
rect 79943 32528 80009 32551
rect 80095 32528 80177 32551
rect 80263 32528 80329 32551
rect 79943 32488 79952 32528
rect 79992 32488 80009 32528
rect 80095 32488 80116 32528
rect 80156 32488 80177 32528
rect 80263 32488 80280 32528
rect 80320 32488 80329 32528
rect 79943 32465 80009 32488
rect 80095 32465 80177 32488
rect 80263 32465 80329 32488
rect 79943 32446 80329 32465
rect 95063 32551 95449 32570
rect 95063 32528 95129 32551
rect 95215 32528 95297 32551
rect 95383 32528 95449 32551
rect 95063 32488 95072 32528
rect 95112 32488 95129 32528
rect 95215 32488 95236 32528
rect 95276 32488 95297 32528
rect 95383 32488 95400 32528
rect 95440 32488 95449 32528
rect 95063 32465 95129 32488
rect 95215 32465 95297 32488
rect 95383 32465 95449 32488
rect 95063 32446 95449 32465
rect 3103 31795 3489 31814
rect 3103 31772 3169 31795
rect 3255 31772 3337 31795
rect 3423 31772 3489 31795
rect 3103 31732 3112 31772
rect 3152 31732 3169 31772
rect 3255 31732 3276 31772
rect 3316 31732 3337 31772
rect 3423 31732 3440 31772
rect 3480 31732 3489 31772
rect 3103 31709 3169 31732
rect 3255 31709 3337 31732
rect 3423 31709 3489 31732
rect 3103 31690 3489 31709
rect 18223 31795 18609 31814
rect 18223 31772 18289 31795
rect 18375 31772 18457 31795
rect 18543 31772 18609 31795
rect 18223 31732 18232 31772
rect 18272 31732 18289 31772
rect 18375 31732 18396 31772
rect 18436 31732 18457 31772
rect 18543 31732 18560 31772
rect 18600 31732 18609 31772
rect 18223 31709 18289 31732
rect 18375 31709 18457 31732
rect 18543 31709 18609 31732
rect 18223 31690 18609 31709
rect 33343 31795 33729 31814
rect 33343 31772 33409 31795
rect 33495 31772 33577 31795
rect 33663 31772 33729 31795
rect 33343 31732 33352 31772
rect 33392 31732 33409 31772
rect 33495 31732 33516 31772
rect 33556 31732 33577 31772
rect 33663 31732 33680 31772
rect 33720 31732 33729 31772
rect 33343 31709 33409 31732
rect 33495 31709 33577 31732
rect 33663 31709 33729 31732
rect 33343 31690 33729 31709
rect 48463 31795 48849 31814
rect 48463 31772 48529 31795
rect 48615 31772 48697 31795
rect 48783 31772 48849 31795
rect 48463 31732 48472 31772
rect 48512 31732 48529 31772
rect 48615 31732 48636 31772
rect 48676 31732 48697 31772
rect 48783 31732 48800 31772
rect 48840 31732 48849 31772
rect 48463 31709 48529 31732
rect 48615 31709 48697 31732
rect 48783 31709 48849 31732
rect 48463 31690 48849 31709
rect 63583 31795 63969 31814
rect 63583 31772 63649 31795
rect 63735 31772 63817 31795
rect 63903 31772 63969 31795
rect 63583 31732 63592 31772
rect 63632 31732 63649 31772
rect 63735 31732 63756 31772
rect 63796 31732 63817 31772
rect 63903 31732 63920 31772
rect 63960 31732 63969 31772
rect 63583 31709 63649 31732
rect 63735 31709 63817 31732
rect 63903 31709 63969 31732
rect 63583 31690 63969 31709
rect 78703 31795 79089 31814
rect 78703 31772 78769 31795
rect 78855 31772 78937 31795
rect 79023 31772 79089 31795
rect 78703 31732 78712 31772
rect 78752 31732 78769 31772
rect 78855 31732 78876 31772
rect 78916 31732 78937 31772
rect 79023 31732 79040 31772
rect 79080 31732 79089 31772
rect 78703 31709 78769 31732
rect 78855 31709 78937 31732
rect 79023 31709 79089 31732
rect 78703 31690 79089 31709
rect 93823 31795 94209 31814
rect 93823 31772 93889 31795
rect 93975 31772 94057 31795
rect 94143 31772 94209 31795
rect 93823 31732 93832 31772
rect 93872 31732 93889 31772
rect 93975 31732 93996 31772
rect 94036 31732 94057 31772
rect 94143 31732 94160 31772
rect 94200 31732 94209 31772
rect 93823 31709 93889 31732
rect 93975 31709 94057 31732
rect 94143 31709 94209 31732
rect 93823 31690 94209 31709
rect 4343 31039 4729 31058
rect 4343 31016 4409 31039
rect 4495 31016 4577 31039
rect 4663 31016 4729 31039
rect 4343 30976 4352 31016
rect 4392 30976 4409 31016
rect 4495 30976 4516 31016
rect 4556 30976 4577 31016
rect 4663 30976 4680 31016
rect 4720 30976 4729 31016
rect 4343 30953 4409 30976
rect 4495 30953 4577 30976
rect 4663 30953 4729 30976
rect 4343 30934 4729 30953
rect 19463 31039 19849 31058
rect 19463 31016 19529 31039
rect 19615 31016 19697 31039
rect 19783 31016 19849 31039
rect 19463 30976 19472 31016
rect 19512 30976 19529 31016
rect 19615 30976 19636 31016
rect 19676 30976 19697 31016
rect 19783 30976 19800 31016
rect 19840 30976 19849 31016
rect 19463 30953 19529 30976
rect 19615 30953 19697 30976
rect 19783 30953 19849 30976
rect 19463 30934 19849 30953
rect 34583 31039 34969 31058
rect 34583 31016 34649 31039
rect 34735 31016 34817 31039
rect 34903 31016 34969 31039
rect 34583 30976 34592 31016
rect 34632 30976 34649 31016
rect 34735 30976 34756 31016
rect 34796 30976 34817 31016
rect 34903 30976 34920 31016
rect 34960 30976 34969 31016
rect 34583 30953 34649 30976
rect 34735 30953 34817 30976
rect 34903 30953 34969 30976
rect 34583 30934 34969 30953
rect 49703 31039 50089 31058
rect 49703 31016 49769 31039
rect 49855 31016 49937 31039
rect 50023 31016 50089 31039
rect 49703 30976 49712 31016
rect 49752 30976 49769 31016
rect 49855 30976 49876 31016
rect 49916 30976 49937 31016
rect 50023 30976 50040 31016
rect 50080 30976 50089 31016
rect 49703 30953 49769 30976
rect 49855 30953 49937 30976
rect 50023 30953 50089 30976
rect 49703 30934 50089 30953
rect 64823 31039 65209 31058
rect 64823 31016 64889 31039
rect 64975 31016 65057 31039
rect 65143 31016 65209 31039
rect 64823 30976 64832 31016
rect 64872 30976 64889 31016
rect 64975 30976 64996 31016
rect 65036 30976 65057 31016
rect 65143 30976 65160 31016
rect 65200 30976 65209 31016
rect 64823 30953 64889 30976
rect 64975 30953 65057 30976
rect 65143 30953 65209 30976
rect 64823 30934 65209 30953
rect 79943 31039 80329 31058
rect 79943 31016 80009 31039
rect 80095 31016 80177 31039
rect 80263 31016 80329 31039
rect 79943 30976 79952 31016
rect 79992 30976 80009 31016
rect 80095 30976 80116 31016
rect 80156 30976 80177 31016
rect 80263 30976 80280 31016
rect 80320 30976 80329 31016
rect 79943 30953 80009 30976
rect 80095 30953 80177 30976
rect 80263 30953 80329 30976
rect 79943 30934 80329 30953
rect 95063 31039 95449 31058
rect 95063 31016 95129 31039
rect 95215 31016 95297 31039
rect 95383 31016 95449 31039
rect 95063 30976 95072 31016
rect 95112 30976 95129 31016
rect 95215 30976 95236 31016
rect 95276 30976 95297 31016
rect 95383 30976 95400 31016
rect 95440 30976 95449 31016
rect 95063 30953 95129 30976
rect 95215 30953 95297 30976
rect 95383 30953 95449 30976
rect 95063 30934 95449 30953
rect 3103 30283 3489 30302
rect 3103 30260 3169 30283
rect 3255 30260 3337 30283
rect 3423 30260 3489 30283
rect 3103 30220 3112 30260
rect 3152 30220 3169 30260
rect 3255 30220 3276 30260
rect 3316 30220 3337 30260
rect 3423 30220 3440 30260
rect 3480 30220 3489 30260
rect 3103 30197 3169 30220
rect 3255 30197 3337 30220
rect 3423 30197 3489 30220
rect 3103 30178 3489 30197
rect 18223 30283 18609 30302
rect 18223 30260 18289 30283
rect 18375 30260 18457 30283
rect 18543 30260 18609 30283
rect 18223 30220 18232 30260
rect 18272 30220 18289 30260
rect 18375 30220 18396 30260
rect 18436 30220 18457 30260
rect 18543 30220 18560 30260
rect 18600 30220 18609 30260
rect 18223 30197 18289 30220
rect 18375 30197 18457 30220
rect 18543 30197 18609 30220
rect 18223 30178 18609 30197
rect 33343 30283 33729 30302
rect 33343 30260 33409 30283
rect 33495 30260 33577 30283
rect 33663 30260 33729 30283
rect 33343 30220 33352 30260
rect 33392 30220 33409 30260
rect 33495 30220 33516 30260
rect 33556 30220 33577 30260
rect 33663 30220 33680 30260
rect 33720 30220 33729 30260
rect 33343 30197 33409 30220
rect 33495 30197 33577 30220
rect 33663 30197 33729 30220
rect 33343 30178 33729 30197
rect 48463 30283 48849 30302
rect 48463 30260 48529 30283
rect 48615 30260 48697 30283
rect 48783 30260 48849 30283
rect 48463 30220 48472 30260
rect 48512 30220 48529 30260
rect 48615 30220 48636 30260
rect 48676 30220 48697 30260
rect 48783 30220 48800 30260
rect 48840 30220 48849 30260
rect 48463 30197 48529 30220
rect 48615 30197 48697 30220
rect 48783 30197 48849 30220
rect 48463 30178 48849 30197
rect 63583 30283 63969 30302
rect 63583 30260 63649 30283
rect 63735 30260 63817 30283
rect 63903 30260 63969 30283
rect 63583 30220 63592 30260
rect 63632 30220 63649 30260
rect 63735 30220 63756 30260
rect 63796 30220 63817 30260
rect 63903 30220 63920 30260
rect 63960 30220 63969 30260
rect 63583 30197 63649 30220
rect 63735 30197 63817 30220
rect 63903 30197 63969 30220
rect 63583 30178 63969 30197
rect 78703 30283 79089 30302
rect 78703 30260 78769 30283
rect 78855 30260 78937 30283
rect 79023 30260 79089 30283
rect 78703 30220 78712 30260
rect 78752 30220 78769 30260
rect 78855 30220 78876 30260
rect 78916 30220 78937 30260
rect 79023 30220 79040 30260
rect 79080 30220 79089 30260
rect 78703 30197 78769 30220
rect 78855 30197 78937 30220
rect 79023 30197 79089 30220
rect 78703 30178 79089 30197
rect 93823 30283 94209 30302
rect 93823 30260 93889 30283
rect 93975 30260 94057 30283
rect 94143 30260 94209 30283
rect 93823 30220 93832 30260
rect 93872 30220 93889 30260
rect 93975 30220 93996 30260
rect 94036 30220 94057 30260
rect 94143 30220 94160 30260
rect 94200 30220 94209 30260
rect 93823 30197 93889 30220
rect 93975 30197 94057 30220
rect 94143 30197 94209 30220
rect 93823 30178 94209 30197
rect 4343 29527 4729 29546
rect 4343 29504 4409 29527
rect 4495 29504 4577 29527
rect 4663 29504 4729 29527
rect 4343 29464 4352 29504
rect 4392 29464 4409 29504
rect 4495 29464 4516 29504
rect 4556 29464 4577 29504
rect 4663 29464 4680 29504
rect 4720 29464 4729 29504
rect 4343 29441 4409 29464
rect 4495 29441 4577 29464
rect 4663 29441 4729 29464
rect 4343 29422 4729 29441
rect 19463 29527 19849 29546
rect 19463 29504 19529 29527
rect 19615 29504 19697 29527
rect 19783 29504 19849 29527
rect 19463 29464 19472 29504
rect 19512 29464 19529 29504
rect 19615 29464 19636 29504
rect 19676 29464 19697 29504
rect 19783 29464 19800 29504
rect 19840 29464 19849 29504
rect 19463 29441 19529 29464
rect 19615 29441 19697 29464
rect 19783 29441 19849 29464
rect 19463 29422 19849 29441
rect 34583 29527 34969 29546
rect 34583 29504 34649 29527
rect 34735 29504 34817 29527
rect 34903 29504 34969 29527
rect 34583 29464 34592 29504
rect 34632 29464 34649 29504
rect 34735 29464 34756 29504
rect 34796 29464 34817 29504
rect 34903 29464 34920 29504
rect 34960 29464 34969 29504
rect 34583 29441 34649 29464
rect 34735 29441 34817 29464
rect 34903 29441 34969 29464
rect 34583 29422 34969 29441
rect 49703 29527 50089 29546
rect 49703 29504 49769 29527
rect 49855 29504 49937 29527
rect 50023 29504 50089 29527
rect 49703 29464 49712 29504
rect 49752 29464 49769 29504
rect 49855 29464 49876 29504
rect 49916 29464 49937 29504
rect 50023 29464 50040 29504
rect 50080 29464 50089 29504
rect 49703 29441 49769 29464
rect 49855 29441 49937 29464
rect 50023 29441 50089 29464
rect 49703 29422 50089 29441
rect 64823 29527 65209 29546
rect 64823 29504 64889 29527
rect 64975 29504 65057 29527
rect 65143 29504 65209 29527
rect 64823 29464 64832 29504
rect 64872 29464 64889 29504
rect 64975 29464 64996 29504
rect 65036 29464 65057 29504
rect 65143 29464 65160 29504
rect 65200 29464 65209 29504
rect 64823 29441 64889 29464
rect 64975 29441 65057 29464
rect 65143 29441 65209 29464
rect 64823 29422 65209 29441
rect 79943 29527 80329 29546
rect 79943 29504 80009 29527
rect 80095 29504 80177 29527
rect 80263 29504 80329 29527
rect 79943 29464 79952 29504
rect 79992 29464 80009 29504
rect 80095 29464 80116 29504
rect 80156 29464 80177 29504
rect 80263 29464 80280 29504
rect 80320 29464 80329 29504
rect 79943 29441 80009 29464
rect 80095 29441 80177 29464
rect 80263 29441 80329 29464
rect 79943 29422 80329 29441
rect 95063 29527 95449 29546
rect 95063 29504 95129 29527
rect 95215 29504 95297 29527
rect 95383 29504 95449 29527
rect 95063 29464 95072 29504
rect 95112 29464 95129 29504
rect 95215 29464 95236 29504
rect 95276 29464 95297 29504
rect 95383 29464 95400 29504
rect 95440 29464 95449 29504
rect 95063 29441 95129 29464
rect 95215 29441 95297 29464
rect 95383 29441 95449 29464
rect 95063 29422 95449 29441
rect 3103 28771 3489 28790
rect 3103 28748 3169 28771
rect 3255 28748 3337 28771
rect 3423 28748 3489 28771
rect 3103 28708 3112 28748
rect 3152 28708 3169 28748
rect 3255 28708 3276 28748
rect 3316 28708 3337 28748
rect 3423 28708 3440 28748
rect 3480 28708 3489 28748
rect 3103 28685 3169 28708
rect 3255 28685 3337 28708
rect 3423 28685 3489 28708
rect 3103 28666 3489 28685
rect 18223 28771 18609 28790
rect 18223 28748 18289 28771
rect 18375 28748 18457 28771
rect 18543 28748 18609 28771
rect 18223 28708 18232 28748
rect 18272 28708 18289 28748
rect 18375 28708 18396 28748
rect 18436 28708 18457 28748
rect 18543 28708 18560 28748
rect 18600 28708 18609 28748
rect 18223 28685 18289 28708
rect 18375 28685 18457 28708
rect 18543 28685 18609 28708
rect 18223 28666 18609 28685
rect 33343 28771 33729 28790
rect 33343 28748 33409 28771
rect 33495 28748 33577 28771
rect 33663 28748 33729 28771
rect 33343 28708 33352 28748
rect 33392 28708 33409 28748
rect 33495 28708 33516 28748
rect 33556 28708 33577 28748
rect 33663 28708 33680 28748
rect 33720 28708 33729 28748
rect 33343 28685 33409 28708
rect 33495 28685 33577 28708
rect 33663 28685 33729 28708
rect 33343 28666 33729 28685
rect 48463 28771 48849 28790
rect 48463 28748 48529 28771
rect 48615 28748 48697 28771
rect 48783 28748 48849 28771
rect 48463 28708 48472 28748
rect 48512 28708 48529 28748
rect 48615 28708 48636 28748
rect 48676 28708 48697 28748
rect 48783 28708 48800 28748
rect 48840 28708 48849 28748
rect 48463 28685 48529 28708
rect 48615 28685 48697 28708
rect 48783 28685 48849 28708
rect 48463 28666 48849 28685
rect 63583 28771 63969 28790
rect 63583 28748 63649 28771
rect 63735 28748 63817 28771
rect 63903 28748 63969 28771
rect 63583 28708 63592 28748
rect 63632 28708 63649 28748
rect 63735 28708 63756 28748
rect 63796 28708 63817 28748
rect 63903 28708 63920 28748
rect 63960 28708 63969 28748
rect 63583 28685 63649 28708
rect 63735 28685 63817 28708
rect 63903 28685 63969 28708
rect 63583 28666 63969 28685
rect 78703 28771 79089 28790
rect 78703 28748 78769 28771
rect 78855 28748 78937 28771
rect 79023 28748 79089 28771
rect 78703 28708 78712 28748
rect 78752 28708 78769 28748
rect 78855 28708 78876 28748
rect 78916 28708 78937 28748
rect 79023 28708 79040 28748
rect 79080 28708 79089 28748
rect 78703 28685 78769 28708
rect 78855 28685 78937 28708
rect 79023 28685 79089 28708
rect 78703 28666 79089 28685
rect 93823 28771 94209 28790
rect 93823 28748 93889 28771
rect 93975 28748 94057 28771
rect 94143 28748 94209 28771
rect 93823 28708 93832 28748
rect 93872 28708 93889 28748
rect 93975 28708 93996 28748
rect 94036 28708 94057 28748
rect 94143 28708 94160 28748
rect 94200 28708 94209 28748
rect 93823 28685 93889 28708
rect 93975 28685 94057 28708
rect 94143 28685 94209 28708
rect 93823 28666 94209 28685
rect 4343 28015 4729 28034
rect 4343 27992 4409 28015
rect 4495 27992 4577 28015
rect 4663 27992 4729 28015
rect 4343 27952 4352 27992
rect 4392 27952 4409 27992
rect 4495 27952 4516 27992
rect 4556 27952 4577 27992
rect 4663 27952 4680 27992
rect 4720 27952 4729 27992
rect 4343 27929 4409 27952
rect 4495 27929 4577 27952
rect 4663 27929 4729 27952
rect 4343 27910 4729 27929
rect 19463 28015 19849 28034
rect 19463 27992 19529 28015
rect 19615 27992 19697 28015
rect 19783 27992 19849 28015
rect 19463 27952 19472 27992
rect 19512 27952 19529 27992
rect 19615 27952 19636 27992
rect 19676 27952 19697 27992
rect 19783 27952 19800 27992
rect 19840 27952 19849 27992
rect 19463 27929 19529 27952
rect 19615 27929 19697 27952
rect 19783 27929 19849 27952
rect 19463 27910 19849 27929
rect 34583 28015 34969 28034
rect 34583 27992 34649 28015
rect 34735 27992 34817 28015
rect 34903 27992 34969 28015
rect 34583 27952 34592 27992
rect 34632 27952 34649 27992
rect 34735 27952 34756 27992
rect 34796 27952 34817 27992
rect 34903 27952 34920 27992
rect 34960 27952 34969 27992
rect 34583 27929 34649 27952
rect 34735 27929 34817 27952
rect 34903 27929 34969 27952
rect 34583 27910 34969 27929
rect 49703 28015 50089 28034
rect 49703 27992 49769 28015
rect 49855 27992 49937 28015
rect 50023 27992 50089 28015
rect 49703 27952 49712 27992
rect 49752 27952 49769 27992
rect 49855 27952 49876 27992
rect 49916 27952 49937 27992
rect 50023 27952 50040 27992
rect 50080 27952 50089 27992
rect 49703 27929 49769 27952
rect 49855 27929 49937 27952
rect 50023 27929 50089 27952
rect 49703 27910 50089 27929
rect 64823 28015 65209 28034
rect 64823 27992 64889 28015
rect 64975 27992 65057 28015
rect 65143 27992 65209 28015
rect 64823 27952 64832 27992
rect 64872 27952 64889 27992
rect 64975 27952 64996 27992
rect 65036 27952 65057 27992
rect 65143 27952 65160 27992
rect 65200 27952 65209 27992
rect 64823 27929 64889 27952
rect 64975 27929 65057 27952
rect 65143 27929 65209 27952
rect 64823 27910 65209 27929
rect 79943 28015 80329 28034
rect 79943 27992 80009 28015
rect 80095 27992 80177 28015
rect 80263 27992 80329 28015
rect 79943 27952 79952 27992
rect 79992 27952 80009 27992
rect 80095 27952 80116 27992
rect 80156 27952 80177 27992
rect 80263 27952 80280 27992
rect 80320 27952 80329 27992
rect 79943 27929 80009 27952
rect 80095 27929 80177 27952
rect 80263 27929 80329 27952
rect 79943 27910 80329 27929
rect 95063 28015 95449 28034
rect 95063 27992 95129 28015
rect 95215 27992 95297 28015
rect 95383 27992 95449 28015
rect 95063 27952 95072 27992
rect 95112 27952 95129 27992
rect 95215 27952 95236 27992
rect 95276 27952 95297 27992
rect 95383 27952 95400 27992
rect 95440 27952 95449 27992
rect 95063 27929 95129 27952
rect 95215 27929 95297 27952
rect 95383 27929 95449 27952
rect 95063 27910 95449 27929
rect 3103 27259 3489 27278
rect 3103 27236 3169 27259
rect 3255 27236 3337 27259
rect 3423 27236 3489 27259
rect 3103 27196 3112 27236
rect 3152 27196 3169 27236
rect 3255 27196 3276 27236
rect 3316 27196 3337 27236
rect 3423 27196 3440 27236
rect 3480 27196 3489 27236
rect 3103 27173 3169 27196
rect 3255 27173 3337 27196
rect 3423 27173 3489 27196
rect 3103 27154 3489 27173
rect 18223 27259 18609 27278
rect 18223 27236 18289 27259
rect 18375 27236 18457 27259
rect 18543 27236 18609 27259
rect 18223 27196 18232 27236
rect 18272 27196 18289 27236
rect 18375 27196 18396 27236
rect 18436 27196 18457 27236
rect 18543 27196 18560 27236
rect 18600 27196 18609 27236
rect 18223 27173 18289 27196
rect 18375 27173 18457 27196
rect 18543 27173 18609 27196
rect 18223 27154 18609 27173
rect 33343 27259 33729 27278
rect 33343 27236 33409 27259
rect 33495 27236 33577 27259
rect 33663 27236 33729 27259
rect 33343 27196 33352 27236
rect 33392 27196 33409 27236
rect 33495 27196 33516 27236
rect 33556 27196 33577 27236
rect 33663 27196 33680 27236
rect 33720 27196 33729 27236
rect 33343 27173 33409 27196
rect 33495 27173 33577 27196
rect 33663 27173 33729 27196
rect 33343 27154 33729 27173
rect 48463 27259 48849 27278
rect 48463 27236 48529 27259
rect 48615 27236 48697 27259
rect 48783 27236 48849 27259
rect 48463 27196 48472 27236
rect 48512 27196 48529 27236
rect 48615 27196 48636 27236
rect 48676 27196 48697 27236
rect 48783 27196 48800 27236
rect 48840 27196 48849 27236
rect 48463 27173 48529 27196
rect 48615 27173 48697 27196
rect 48783 27173 48849 27196
rect 48463 27154 48849 27173
rect 63583 27259 63969 27278
rect 63583 27236 63649 27259
rect 63735 27236 63817 27259
rect 63903 27236 63969 27259
rect 63583 27196 63592 27236
rect 63632 27196 63649 27236
rect 63735 27196 63756 27236
rect 63796 27196 63817 27236
rect 63903 27196 63920 27236
rect 63960 27196 63969 27236
rect 63583 27173 63649 27196
rect 63735 27173 63817 27196
rect 63903 27173 63969 27196
rect 63583 27154 63969 27173
rect 78703 27259 79089 27278
rect 78703 27236 78769 27259
rect 78855 27236 78937 27259
rect 79023 27236 79089 27259
rect 78703 27196 78712 27236
rect 78752 27196 78769 27236
rect 78855 27196 78876 27236
rect 78916 27196 78937 27236
rect 79023 27196 79040 27236
rect 79080 27196 79089 27236
rect 78703 27173 78769 27196
rect 78855 27173 78937 27196
rect 79023 27173 79089 27196
rect 78703 27154 79089 27173
rect 93823 27259 94209 27278
rect 93823 27236 93889 27259
rect 93975 27236 94057 27259
rect 94143 27236 94209 27259
rect 93823 27196 93832 27236
rect 93872 27196 93889 27236
rect 93975 27196 93996 27236
rect 94036 27196 94057 27236
rect 94143 27196 94160 27236
rect 94200 27196 94209 27236
rect 93823 27173 93889 27196
rect 93975 27173 94057 27196
rect 94143 27173 94209 27196
rect 93823 27154 94209 27173
rect 4343 26503 4729 26522
rect 4343 26480 4409 26503
rect 4495 26480 4577 26503
rect 4663 26480 4729 26503
rect 4343 26440 4352 26480
rect 4392 26440 4409 26480
rect 4495 26440 4516 26480
rect 4556 26440 4577 26480
rect 4663 26440 4680 26480
rect 4720 26440 4729 26480
rect 4343 26417 4409 26440
rect 4495 26417 4577 26440
rect 4663 26417 4729 26440
rect 4343 26398 4729 26417
rect 19463 26503 19849 26522
rect 19463 26480 19529 26503
rect 19615 26480 19697 26503
rect 19783 26480 19849 26503
rect 19463 26440 19472 26480
rect 19512 26440 19529 26480
rect 19615 26440 19636 26480
rect 19676 26440 19697 26480
rect 19783 26440 19800 26480
rect 19840 26440 19849 26480
rect 19463 26417 19529 26440
rect 19615 26417 19697 26440
rect 19783 26417 19849 26440
rect 19463 26398 19849 26417
rect 34583 26503 34969 26522
rect 34583 26480 34649 26503
rect 34735 26480 34817 26503
rect 34903 26480 34969 26503
rect 34583 26440 34592 26480
rect 34632 26440 34649 26480
rect 34735 26440 34756 26480
rect 34796 26440 34817 26480
rect 34903 26440 34920 26480
rect 34960 26440 34969 26480
rect 34583 26417 34649 26440
rect 34735 26417 34817 26440
rect 34903 26417 34969 26440
rect 34583 26398 34969 26417
rect 49703 26503 50089 26522
rect 49703 26480 49769 26503
rect 49855 26480 49937 26503
rect 50023 26480 50089 26503
rect 49703 26440 49712 26480
rect 49752 26440 49769 26480
rect 49855 26440 49876 26480
rect 49916 26440 49937 26480
rect 50023 26440 50040 26480
rect 50080 26440 50089 26480
rect 49703 26417 49769 26440
rect 49855 26417 49937 26440
rect 50023 26417 50089 26440
rect 49703 26398 50089 26417
rect 64823 26503 65209 26522
rect 64823 26480 64889 26503
rect 64975 26480 65057 26503
rect 65143 26480 65209 26503
rect 64823 26440 64832 26480
rect 64872 26440 64889 26480
rect 64975 26440 64996 26480
rect 65036 26440 65057 26480
rect 65143 26440 65160 26480
rect 65200 26440 65209 26480
rect 64823 26417 64889 26440
rect 64975 26417 65057 26440
rect 65143 26417 65209 26440
rect 64823 26398 65209 26417
rect 79943 26503 80329 26522
rect 79943 26480 80009 26503
rect 80095 26480 80177 26503
rect 80263 26480 80329 26503
rect 79943 26440 79952 26480
rect 79992 26440 80009 26480
rect 80095 26440 80116 26480
rect 80156 26440 80177 26480
rect 80263 26440 80280 26480
rect 80320 26440 80329 26480
rect 79943 26417 80009 26440
rect 80095 26417 80177 26440
rect 80263 26417 80329 26440
rect 79943 26398 80329 26417
rect 95063 26503 95449 26522
rect 95063 26480 95129 26503
rect 95215 26480 95297 26503
rect 95383 26480 95449 26503
rect 95063 26440 95072 26480
rect 95112 26440 95129 26480
rect 95215 26440 95236 26480
rect 95276 26440 95297 26480
rect 95383 26440 95400 26480
rect 95440 26440 95449 26480
rect 95063 26417 95129 26440
rect 95215 26417 95297 26440
rect 95383 26417 95449 26440
rect 95063 26398 95449 26417
rect 3103 25747 3489 25766
rect 3103 25724 3169 25747
rect 3255 25724 3337 25747
rect 3423 25724 3489 25747
rect 3103 25684 3112 25724
rect 3152 25684 3169 25724
rect 3255 25684 3276 25724
rect 3316 25684 3337 25724
rect 3423 25684 3440 25724
rect 3480 25684 3489 25724
rect 3103 25661 3169 25684
rect 3255 25661 3337 25684
rect 3423 25661 3489 25684
rect 3103 25642 3489 25661
rect 18223 25747 18609 25766
rect 18223 25724 18289 25747
rect 18375 25724 18457 25747
rect 18543 25724 18609 25747
rect 18223 25684 18232 25724
rect 18272 25684 18289 25724
rect 18375 25684 18396 25724
rect 18436 25684 18457 25724
rect 18543 25684 18560 25724
rect 18600 25684 18609 25724
rect 18223 25661 18289 25684
rect 18375 25661 18457 25684
rect 18543 25661 18609 25684
rect 18223 25642 18609 25661
rect 33343 25747 33729 25766
rect 33343 25724 33409 25747
rect 33495 25724 33577 25747
rect 33663 25724 33729 25747
rect 33343 25684 33352 25724
rect 33392 25684 33409 25724
rect 33495 25684 33516 25724
rect 33556 25684 33577 25724
rect 33663 25684 33680 25724
rect 33720 25684 33729 25724
rect 33343 25661 33409 25684
rect 33495 25661 33577 25684
rect 33663 25661 33729 25684
rect 33343 25642 33729 25661
rect 48463 25747 48849 25766
rect 48463 25724 48529 25747
rect 48615 25724 48697 25747
rect 48783 25724 48849 25747
rect 48463 25684 48472 25724
rect 48512 25684 48529 25724
rect 48615 25684 48636 25724
rect 48676 25684 48697 25724
rect 48783 25684 48800 25724
rect 48840 25684 48849 25724
rect 48463 25661 48529 25684
rect 48615 25661 48697 25684
rect 48783 25661 48849 25684
rect 48463 25642 48849 25661
rect 63583 25747 63969 25766
rect 63583 25724 63649 25747
rect 63735 25724 63817 25747
rect 63903 25724 63969 25747
rect 63583 25684 63592 25724
rect 63632 25684 63649 25724
rect 63735 25684 63756 25724
rect 63796 25684 63817 25724
rect 63903 25684 63920 25724
rect 63960 25684 63969 25724
rect 63583 25661 63649 25684
rect 63735 25661 63817 25684
rect 63903 25661 63969 25684
rect 63583 25642 63969 25661
rect 78703 25747 79089 25766
rect 78703 25724 78769 25747
rect 78855 25724 78937 25747
rect 79023 25724 79089 25747
rect 78703 25684 78712 25724
rect 78752 25684 78769 25724
rect 78855 25684 78876 25724
rect 78916 25684 78937 25724
rect 79023 25684 79040 25724
rect 79080 25684 79089 25724
rect 78703 25661 78769 25684
rect 78855 25661 78937 25684
rect 79023 25661 79089 25684
rect 78703 25642 79089 25661
rect 93823 25747 94209 25766
rect 93823 25724 93889 25747
rect 93975 25724 94057 25747
rect 94143 25724 94209 25747
rect 93823 25684 93832 25724
rect 93872 25684 93889 25724
rect 93975 25684 93996 25724
rect 94036 25684 94057 25724
rect 94143 25684 94160 25724
rect 94200 25684 94209 25724
rect 93823 25661 93889 25684
rect 93975 25661 94057 25684
rect 94143 25661 94209 25684
rect 93823 25642 94209 25661
rect 4343 24991 4729 25010
rect 4343 24968 4409 24991
rect 4495 24968 4577 24991
rect 4663 24968 4729 24991
rect 4343 24928 4352 24968
rect 4392 24928 4409 24968
rect 4495 24928 4516 24968
rect 4556 24928 4577 24968
rect 4663 24928 4680 24968
rect 4720 24928 4729 24968
rect 4343 24905 4409 24928
rect 4495 24905 4577 24928
rect 4663 24905 4729 24928
rect 4343 24886 4729 24905
rect 19463 24991 19849 25010
rect 19463 24968 19529 24991
rect 19615 24968 19697 24991
rect 19783 24968 19849 24991
rect 19463 24928 19472 24968
rect 19512 24928 19529 24968
rect 19615 24928 19636 24968
rect 19676 24928 19697 24968
rect 19783 24928 19800 24968
rect 19840 24928 19849 24968
rect 19463 24905 19529 24928
rect 19615 24905 19697 24928
rect 19783 24905 19849 24928
rect 19463 24886 19849 24905
rect 34583 24991 34969 25010
rect 34583 24968 34649 24991
rect 34735 24968 34817 24991
rect 34903 24968 34969 24991
rect 34583 24928 34592 24968
rect 34632 24928 34649 24968
rect 34735 24928 34756 24968
rect 34796 24928 34817 24968
rect 34903 24928 34920 24968
rect 34960 24928 34969 24968
rect 34583 24905 34649 24928
rect 34735 24905 34817 24928
rect 34903 24905 34969 24928
rect 34583 24886 34969 24905
rect 49703 24991 50089 25010
rect 49703 24968 49769 24991
rect 49855 24968 49937 24991
rect 50023 24968 50089 24991
rect 49703 24928 49712 24968
rect 49752 24928 49769 24968
rect 49855 24928 49876 24968
rect 49916 24928 49937 24968
rect 50023 24928 50040 24968
rect 50080 24928 50089 24968
rect 49703 24905 49769 24928
rect 49855 24905 49937 24928
rect 50023 24905 50089 24928
rect 49703 24886 50089 24905
rect 64823 24991 65209 25010
rect 64823 24968 64889 24991
rect 64975 24968 65057 24991
rect 65143 24968 65209 24991
rect 64823 24928 64832 24968
rect 64872 24928 64889 24968
rect 64975 24928 64996 24968
rect 65036 24928 65057 24968
rect 65143 24928 65160 24968
rect 65200 24928 65209 24968
rect 64823 24905 64889 24928
rect 64975 24905 65057 24928
rect 65143 24905 65209 24928
rect 64823 24886 65209 24905
rect 79943 24991 80329 25010
rect 79943 24968 80009 24991
rect 80095 24968 80177 24991
rect 80263 24968 80329 24991
rect 79943 24928 79952 24968
rect 79992 24928 80009 24968
rect 80095 24928 80116 24968
rect 80156 24928 80177 24968
rect 80263 24928 80280 24968
rect 80320 24928 80329 24968
rect 79943 24905 80009 24928
rect 80095 24905 80177 24928
rect 80263 24905 80329 24928
rect 79943 24886 80329 24905
rect 95063 24991 95449 25010
rect 95063 24968 95129 24991
rect 95215 24968 95297 24991
rect 95383 24968 95449 24991
rect 95063 24928 95072 24968
rect 95112 24928 95129 24968
rect 95215 24928 95236 24968
rect 95276 24928 95297 24968
rect 95383 24928 95400 24968
rect 95440 24928 95449 24968
rect 95063 24905 95129 24928
rect 95215 24905 95297 24928
rect 95383 24905 95449 24928
rect 95063 24886 95449 24905
rect 3103 24235 3489 24254
rect 3103 24212 3169 24235
rect 3255 24212 3337 24235
rect 3423 24212 3489 24235
rect 3103 24172 3112 24212
rect 3152 24172 3169 24212
rect 3255 24172 3276 24212
rect 3316 24172 3337 24212
rect 3423 24172 3440 24212
rect 3480 24172 3489 24212
rect 3103 24149 3169 24172
rect 3255 24149 3337 24172
rect 3423 24149 3489 24172
rect 3103 24130 3489 24149
rect 18223 24235 18609 24254
rect 18223 24212 18289 24235
rect 18375 24212 18457 24235
rect 18543 24212 18609 24235
rect 18223 24172 18232 24212
rect 18272 24172 18289 24212
rect 18375 24172 18396 24212
rect 18436 24172 18457 24212
rect 18543 24172 18560 24212
rect 18600 24172 18609 24212
rect 18223 24149 18289 24172
rect 18375 24149 18457 24172
rect 18543 24149 18609 24172
rect 18223 24130 18609 24149
rect 33343 24235 33729 24254
rect 33343 24212 33409 24235
rect 33495 24212 33577 24235
rect 33663 24212 33729 24235
rect 33343 24172 33352 24212
rect 33392 24172 33409 24212
rect 33495 24172 33516 24212
rect 33556 24172 33577 24212
rect 33663 24172 33680 24212
rect 33720 24172 33729 24212
rect 33343 24149 33409 24172
rect 33495 24149 33577 24172
rect 33663 24149 33729 24172
rect 33343 24130 33729 24149
rect 48463 24235 48849 24254
rect 48463 24212 48529 24235
rect 48615 24212 48697 24235
rect 48783 24212 48849 24235
rect 48463 24172 48472 24212
rect 48512 24172 48529 24212
rect 48615 24172 48636 24212
rect 48676 24172 48697 24212
rect 48783 24172 48800 24212
rect 48840 24172 48849 24212
rect 48463 24149 48529 24172
rect 48615 24149 48697 24172
rect 48783 24149 48849 24172
rect 48463 24130 48849 24149
rect 63583 24235 63969 24254
rect 63583 24212 63649 24235
rect 63735 24212 63817 24235
rect 63903 24212 63969 24235
rect 63583 24172 63592 24212
rect 63632 24172 63649 24212
rect 63735 24172 63756 24212
rect 63796 24172 63817 24212
rect 63903 24172 63920 24212
rect 63960 24172 63969 24212
rect 63583 24149 63649 24172
rect 63735 24149 63817 24172
rect 63903 24149 63969 24172
rect 63583 24130 63969 24149
rect 78703 24235 79089 24254
rect 78703 24212 78769 24235
rect 78855 24212 78937 24235
rect 79023 24212 79089 24235
rect 78703 24172 78712 24212
rect 78752 24172 78769 24212
rect 78855 24172 78876 24212
rect 78916 24172 78937 24212
rect 79023 24172 79040 24212
rect 79080 24172 79089 24212
rect 78703 24149 78769 24172
rect 78855 24149 78937 24172
rect 79023 24149 79089 24172
rect 78703 24130 79089 24149
rect 93823 24235 94209 24254
rect 93823 24212 93889 24235
rect 93975 24212 94057 24235
rect 94143 24212 94209 24235
rect 93823 24172 93832 24212
rect 93872 24172 93889 24212
rect 93975 24172 93996 24212
rect 94036 24172 94057 24212
rect 94143 24172 94160 24212
rect 94200 24172 94209 24212
rect 93823 24149 93889 24172
rect 93975 24149 94057 24172
rect 94143 24149 94209 24172
rect 93823 24130 94209 24149
rect 4343 23479 4729 23498
rect 4343 23456 4409 23479
rect 4495 23456 4577 23479
rect 4663 23456 4729 23479
rect 4343 23416 4352 23456
rect 4392 23416 4409 23456
rect 4495 23416 4516 23456
rect 4556 23416 4577 23456
rect 4663 23416 4680 23456
rect 4720 23416 4729 23456
rect 4343 23393 4409 23416
rect 4495 23393 4577 23416
rect 4663 23393 4729 23416
rect 4343 23374 4729 23393
rect 19463 23479 19849 23498
rect 19463 23456 19529 23479
rect 19615 23456 19697 23479
rect 19783 23456 19849 23479
rect 19463 23416 19472 23456
rect 19512 23416 19529 23456
rect 19615 23416 19636 23456
rect 19676 23416 19697 23456
rect 19783 23416 19800 23456
rect 19840 23416 19849 23456
rect 19463 23393 19529 23416
rect 19615 23393 19697 23416
rect 19783 23393 19849 23416
rect 19463 23374 19849 23393
rect 34583 23479 34969 23498
rect 34583 23456 34649 23479
rect 34735 23456 34817 23479
rect 34903 23456 34969 23479
rect 34583 23416 34592 23456
rect 34632 23416 34649 23456
rect 34735 23416 34756 23456
rect 34796 23416 34817 23456
rect 34903 23416 34920 23456
rect 34960 23416 34969 23456
rect 34583 23393 34649 23416
rect 34735 23393 34817 23416
rect 34903 23393 34969 23416
rect 34583 23374 34969 23393
rect 49703 23479 50089 23498
rect 49703 23456 49769 23479
rect 49855 23456 49937 23479
rect 50023 23456 50089 23479
rect 49703 23416 49712 23456
rect 49752 23416 49769 23456
rect 49855 23416 49876 23456
rect 49916 23416 49937 23456
rect 50023 23416 50040 23456
rect 50080 23416 50089 23456
rect 49703 23393 49769 23416
rect 49855 23393 49937 23416
rect 50023 23393 50089 23416
rect 49703 23374 50089 23393
rect 64823 23479 65209 23498
rect 64823 23456 64889 23479
rect 64975 23456 65057 23479
rect 65143 23456 65209 23479
rect 64823 23416 64832 23456
rect 64872 23416 64889 23456
rect 64975 23416 64996 23456
rect 65036 23416 65057 23456
rect 65143 23416 65160 23456
rect 65200 23416 65209 23456
rect 64823 23393 64889 23416
rect 64975 23393 65057 23416
rect 65143 23393 65209 23416
rect 64823 23374 65209 23393
rect 79943 23479 80329 23498
rect 79943 23456 80009 23479
rect 80095 23456 80177 23479
rect 80263 23456 80329 23479
rect 79943 23416 79952 23456
rect 79992 23416 80009 23456
rect 80095 23416 80116 23456
rect 80156 23416 80177 23456
rect 80263 23416 80280 23456
rect 80320 23416 80329 23456
rect 79943 23393 80009 23416
rect 80095 23393 80177 23416
rect 80263 23393 80329 23416
rect 79943 23374 80329 23393
rect 95063 23479 95449 23498
rect 95063 23456 95129 23479
rect 95215 23456 95297 23479
rect 95383 23456 95449 23479
rect 95063 23416 95072 23456
rect 95112 23416 95129 23456
rect 95215 23416 95236 23456
rect 95276 23416 95297 23456
rect 95383 23416 95400 23456
rect 95440 23416 95449 23456
rect 95063 23393 95129 23416
rect 95215 23393 95297 23416
rect 95383 23393 95449 23416
rect 95063 23374 95449 23393
rect 3103 22723 3489 22742
rect 3103 22700 3169 22723
rect 3255 22700 3337 22723
rect 3423 22700 3489 22723
rect 3103 22660 3112 22700
rect 3152 22660 3169 22700
rect 3255 22660 3276 22700
rect 3316 22660 3337 22700
rect 3423 22660 3440 22700
rect 3480 22660 3489 22700
rect 3103 22637 3169 22660
rect 3255 22637 3337 22660
rect 3423 22637 3489 22660
rect 3103 22618 3489 22637
rect 18223 22723 18609 22742
rect 18223 22700 18289 22723
rect 18375 22700 18457 22723
rect 18543 22700 18609 22723
rect 18223 22660 18232 22700
rect 18272 22660 18289 22700
rect 18375 22660 18396 22700
rect 18436 22660 18457 22700
rect 18543 22660 18560 22700
rect 18600 22660 18609 22700
rect 18223 22637 18289 22660
rect 18375 22637 18457 22660
rect 18543 22637 18609 22660
rect 18223 22618 18609 22637
rect 33343 22723 33729 22742
rect 33343 22700 33409 22723
rect 33495 22700 33577 22723
rect 33663 22700 33729 22723
rect 33343 22660 33352 22700
rect 33392 22660 33409 22700
rect 33495 22660 33516 22700
rect 33556 22660 33577 22700
rect 33663 22660 33680 22700
rect 33720 22660 33729 22700
rect 33343 22637 33409 22660
rect 33495 22637 33577 22660
rect 33663 22637 33729 22660
rect 33343 22618 33729 22637
rect 48463 22723 48849 22742
rect 48463 22700 48529 22723
rect 48615 22700 48697 22723
rect 48783 22700 48849 22723
rect 48463 22660 48472 22700
rect 48512 22660 48529 22700
rect 48615 22660 48636 22700
rect 48676 22660 48697 22700
rect 48783 22660 48800 22700
rect 48840 22660 48849 22700
rect 48463 22637 48529 22660
rect 48615 22637 48697 22660
rect 48783 22637 48849 22660
rect 48463 22618 48849 22637
rect 63583 22723 63969 22742
rect 63583 22700 63649 22723
rect 63735 22700 63817 22723
rect 63903 22700 63969 22723
rect 63583 22660 63592 22700
rect 63632 22660 63649 22700
rect 63735 22660 63756 22700
rect 63796 22660 63817 22700
rect 63903 22660 63920 22700
rect 63960 22660 63969 22700
rect 63583 22637 63649 22660
rect 63735 22637 63817 22660
rect 63903 22637 63969 22660
rect 63583 22618 63969 22637
rect 78703 22723 79089 22742
rect 78703 22700 78769 22723
rect 78855 22700 78937 22723
rect 79023 22700 79089 22723
rect 78703 22660 78712 22700
rect 78752 22660 78769 22700
rect 78855 22660 78876 22700
rect 78916 22660 78937 22700
rect 79023 22660 79040 22700
rect 79080 22660 79089 22700
rect 78703 22637 78769 22660
rect 78855 22637 78937 22660
rect 79023 22637 79089 22660
rect 78703 22618 79089 22637
rect 93823 22723 94209 22742
rect 93823 22700 93889 22723
rect 93975 22700 94057 22723
rect 94143 22700 94209 22723
rect 93823 22660 93832 22700
rect 93872 22660 93889 22700
rect 93975 22660 93996 22700
rect 94036 22660 94057 22700
rect 94143 22660 94160 22700
rect 94200 22660 94209 22700
rect 93823 22637 93889 22660
rect 93975 22637 94057 22660
rect 94143 22637 94209 22660
rect 93823 22618 94209 22637
rect 4343 21967 4729 21986
rect 4343 21944 4409 21967
rect 4495 21944 4577 21967
rect 4663 21944 4729 21967
rect 4343 21904 4352 21944
rect 4392 21904 4409 21944
rect 4495 21904 4516 21944
rect 4556 21904 4577 21944
rect 4663 21904 4680 21944
rect 4720 21904 4729 21944
rect 4343 21881 4409 21904
rect 4495 21881 4577 21904
rect 4663 21881 4729 21904
rect 4343 21862 4729 21881
rect 19463 21967 19849 21986
rect 19463 21944 19529 21967
rect 19615 21944 19697 21967
rect 19783 21944 19849 21967
rect 19463 21904 19472 21944
rect 19512 21904 19529 21944
rect 19615 21904 19636 21944
rect 19676 21904 19697 21944
rect 19783 21904 19800 21944
rect 19840 21904 19849 21944
rect 19463 21881 19529 21904
rect 19615 21881 19697 21904
rect 19783 21881 19849 21904
rect 19463 21862 19849 21881
rect 34583 21967 34969 21986
rect 34583 21944 34649 21967
rect 34735 21944 34817 21967
rect 34903 21944 34969 21967
rect 34583 21904 34592 21944
rect 34632 21904 34649 21944
rect 34735 21904 34756 21944
rect 34796 21904 34817 21944
rect 34903 21904 34920 21944
rect 34960 21904 34969 21944
rect 34583 21881 34649 21904
rect 34735 21881 34817 21904
rect 34903 21881 34969 21904
rect 34583 21862 34969 21881
rect 49703 21967 50089 21986
rect 49703 21944 49769 21967
rect 49855 21944 49937 21967
rect 50023 21944 50089 21967
rect 49703 21904 49712 21944
rect 49752 21904 49769 21944
rect 49855 21904 49876 21944
rect 49916 21904 49937 21944
rect 50023 21904 50040 21944
rect 50080 21904 50089 21944
rect 49703 21881 49769 21904
rect 49855 21881 49937 21904
rect 50023 21881 50089 21904
rect 49703 21862 50089 21881
rect 64823 21967 65209 21986
rect 64823 21944 64889 21967
rect 64975 21944 65057 21967
rect 65143 21944 65209 21967
rect 64823 21904 64832 21944
rect 64872 21904 64889 21944
rect 64975 21904 64996 21944
rect 65036 21904 65057 21944
rect 65143 21904 65160 21944
rect 65200 21904 65209 21944
rect 64823 21881 64889 21904
rect 64975 21881 65057 21904
rect 65143 21881 65209 21904
rect 64823 21862 65209 21881
rect 79943 21967 80329 21986
rect 79943 21944 80009 21967
rect 80095 21944 80177 21967
rect 80263 21944 80329 21967
rect 79943 21904 79952 21944
rect 79992 21904 80009 21944
rect 80095 21904 80116 21944
rect 80156 21904 80177 21944
rect 80263 21904 80280 21944
rect 80320 21904 80329 21944
rect 79943 21881 80009 21904
rect 80095 21881 80177 21904
rect 80263 21881 80329 21904
rect 79943 21862 80329 21881
rect 95063 21967 95449 21986
rect 95063 21944 95129 21967
rect 95215 21944 95297 21967
rect 95383 21944 95449 21967
rect 95063 21904 95072 21944
rect 95112 21904 95129 21944
rect 95215 21904 95236 21944
rect 95276 21904 95297 21944
rect 95383 21904 95400 21944
rect 95440 21904 95449 21944
rect 95063 21881 95129 21904
rect 95215 21881 95297 21904
rect 95383 21881 95449 21904
rect 95063 21862 95449 21881
rect 3103 21211 3489 21230
rect 3103 21188 3169 21211
rect 3255 21188 3337 21211
rect 3423 21188 3489 21211
rect 3103 21148 3112 21188
rect 3152 21148 3169 21188
rect 3255 21148 3276 21188
rect 3316 21148 3337 21188
rect 3423 21148 3440 21188
rect 3480 21148 3489 21188
rect 3103 21125 3169 21148
rect 3255 21125 3337 21148
rect 3423 21125 3489 21148
rect 3103 21106 3489 21125
rect 18223 21211 18609 21230
rect 18223 21188 18289 21211
rect 18375 21188 18457 21211
rect 18543 21188 18609 21211
rect 18223 21148 18232 21188
rect 18272 21148 18289 21188
rect 18375 21148 18396 21188
rect 18436 21148 18457 21188
rect 18543 21148 18560 21188
rect 18600 21148 18609 21188
rect 18223 21125 18289 21148
rect 18375 21125 18457 21148
rect 18543 21125 18609 21148
rect 18223 21106 18609 21125
rect 33343 21211 33729 21230
rect 33343 21188 33409 21211
rect 33495 21188 33577 21211
rect 33663 21188 33729 21211
rect 33343 21148 33352 21188
rect 33392 21148 33409 21188
rect 33495 21148 33516 21188
rect 33556 21148 33577 21188
rect 33663 21148 33680 21188
rect 33720 21148 33729 21188
rect 33343 21125 33409 21148
rect 33495 21125 33577 21148
rect 33663 21125 33729 21148
rect 33343 21106 33729 21125
rect 48463 21211 48849 21230
rect 48463 21188 48529 21211
rect 48615 21188 48697 21211
rect 48783 21188 48849 21211
rect 48463 21148 48472 21188
rect 48512 21148 48529 21188
rect 48615 21148 48636 21188
rect 48676 21148 48697 21188
rect 48783 21148 48800 21188
rect 48840 21148 48849 21188
rect 48463 21125 48529 21148
rect 48615 21125 48697 21148
rect 48783 21125 48849 21148
rect 48463 21106 48849 21125
rect 63583 21211 63969 21230
rect 63583 21188 63649 21211
rect 63735 21188 63817 21211
rect 63903 21188 63969 21211
rect 63583 21148 63592 21188
rect 63632 21148 63649 21188
rect 63735 21148 63756 21188
rect 63796 21148 63817 21188
rect 63903 21148 63920 21188
rect 63960 21148 63969 21188
rect 63583 21125 63649 21148
rect 63735 21125 63817 21148
rect 63903 21125 63969 21148
rect 63583 21106 63969 21125
rect 78703 21211 79089 21230
rect 78703 21188 78769 21211
rect 78855 21188 78937 21211
rect 79023 21188 79089 21211
rect 78703 21148 78712 21188
rect 78752 21148 78769 21188
rect 78855 21148 78876 21188
rect 78916 21148 78937 21188
rect 79023 21148 79040 21188
rect 79080 21148 79089 21188
rect 78703 21125 78769 21148
rect 78855 21125 78937 21148
rect 79023 21125 79089 21148
rect 78703 21106 79089 21125
rect 93823 21211 94209 21230
rect 93823 21188 93889 21211
rect 93975 21188 94057 21211
rect 94143 21188 94209 21211
rect 93823 21148 93832 21188
rect 93872 21148 93889 21188
rect 93975 21148 93996 21188
rect 94036 21148 94057 21188
rect 94143 21148 94160 21188
rect 94200 21148 94209 21188
rect 93823 21125 93889 21148
rect 93975 21125 94057 21148
rect 94143 21125 94209 21148
rect 93823 21106 94209 21125
rect 4343 20455 4729 20474
rect 4343 20432 4409 20455
rect 4495 20432 4577 20455
rect 4663 20432 4729 20455
rect 4343 20392 4352 20432
rect 4392 20392 4409 20432
rect 4495 20392 4516 20432
rect 4556 20392 4577 20432
rect 4663 20392 4680 20432
rect 4720 20392 4729 20432
rect 4343 20369 4409 20392
rect 4495 20369 4577 20392
rect 4663 20369 4729 20392
rect 4343 20350 4729 20369
rect 19463 20455 19849 20474
rect 19463 20432 19529 20455
rect 19615 20432 19697 20455
rect 19783 20432 19849 20455
rect 19463 20392 19472 20432
rect 19512 20392 19529 20432
rect 19615 20392 19636 20432
rect 19676 20392 19697 20432
rect 19783 20392 19800 20432
rect 19840 20392 19849 20432
rect 19463 20369 19529 20392
rect 19615 20369 19697 20392
rect 19783 20369 19849 20392
rect 19463 20350 19849 20369
rect 34583 20455 34969 20474
rect 34583 20432 34649 20455
rect 34735 20432 34817 20455
rect 34903 20432 34969 20455
rect 34583 20392 34592 20432
rect 34632 20392 34649 20432
rect 34735 20392 34756 20432
rect 34796 20392 34817 20432
rect 34903 20392 34920 20432
rect 34960 20392 34969 20432
rect 34583 20369 34649 20392
rect 34735 20369 34817 20392
rect 34903 20369 34969 20392
rect 34583 20350 34969 20369
rect 49703 20455 50089 20474
rect 49703 20432 49769 20455
rect 49855 20432 49937 20455
rect 50023 20432 50089 20455
rect 49703 20392 49712 20432
rect 49752 20392 49769 20432
rect 49855 20392 49876 20432
rect 49916 20392 49937 20432
rect 50023 20392 50040 20432
rect 50080 20392 50089 20432
rect 49703 20369 49769 20392
rect 49855 20369 49937 20392
rect 50023 20369 50089 20392
rect 49703 20350 50089 20369
rect 64823 20455 65209 20474
rect 64823 20432 64889 20455
rect 64975 20432 65057 20455
rect 65143 20432 65209 20455
rect 64823 20392 64832 20432
rect 64872 20392 64889 20432
rect 64975 20392 64996 20432
rect 65036 20392 65057 20432
rect 65143 20392 65160 20432
rect 65200 20392 65209 20432
rect 64823 20369 64889 20392
rect 64975 20369 65057 20392
rect 65143 20369 65209 20392
rect 64823 20350 65209 20369
rect 79943 20455 80329 20474
rect 79943 20432 80009 20455
rect 80095 20432 80177 20455
rect 80263 20432 80329 20455
rect 79943 20392 79952 20432
rect 79992 20392 80009 20432
rect 80095 20392 80116 20432
rect 80156 20392 80177 20432
rect 80263 20392 80280 20432
rect 80320 20392 80329 20432
rect 79943 20369 80009 20392
rect 80095 20369 80177 20392
rect 80263 20369 80329 20392
rect 79943 20350 80329 20369
rect 95063 20455 95449 20474
rect 95063 20432 95129 20455
rect 95215 20432 95297 20455
rect 95383 20432 95449 20455
rect 95063 20392 95072 20432
rect 95112 20392 95129 20432
rect 95215 20392 95236 20432
rect 95276 20392 95297 20432
rect 95383 20392 95400 20432
rect 95440 20392 95449 20432
rect 95063 20369 95129 20392
rect 95215 20369 95297 20392
rect 95383 20369 95449 20392
rect 95063 20350 95449 20369
rect 3103 19699 3489 19718
rect 3103 19676 3169 19699
rect 3255 19676 3337 19699
rect 3423 19676 3489 19699
rect 3103 19636 3112 19676
rect 3152 19636 3169 19676
rect 3255 19636 3276 19676
rect 3316 19636 3337 19676
rect 3423 19636 3440 19676
rect 3480 19636 3489 19676
rect 3103 19613 3169 19636
rect 3255 19613 3337 19636
rect 3423 19613 3489 19636
rect 3103 19594 3489 19613
rect 18223 19699 18609 19718
rect 18223 19676 18289 19699
rect 18375 19676 18457 19699
rect 18543 19676 18609 19699
rect 18223 19636 18232 19676
rect 18272 19636 18289 19676
rect 18375 19636 18396 19676
rect 18436 19636 18457 19676
rect 18543 19636 18560 19676
rect 18600 19636 18609 19676
rect 18223 19613 18289 19636
rect 18375 19613 18457 19636
rect 18543 19613 18609 19636
rect 18223 19594 18609 19613
rect 33343 19699 33729 19718
rect 33343 19676 33409 19699
rect 33495 19676 33577 19699
rect 33663 19676 33729 19699
rect 33343 19636 33352 19676
rect 33392 19636 33409 19676
rect 33495 19636 33516 19676
rect 33556 19636 33577 19676
rect 33663 19636 33680 19676
rect 33720 19636 33729 19676
rect 33343 19613 33409 19636
rect 33495 19613 33577 19636
rect 33663 19613 33729 19636
rect 33343 19594 33729 19613
rect 48463 19699 48849 19718
rect 48463 19676 48529 19699
rect 48615 19676 48697 19699
rect 48783 19676 48849 19699
rect 48463 19636 48472 19676
rect 48512 19636 48529 19676
rect 48615 19636 48636 19676
rect 48676 19636 48697 19676
rect 48783 19636 48800 19676
rect 48840 19636 48849 19676
rect 48463 19613 48529 19636
rect 48615 19613 48697 19636
rect 48783 19613 48849 19636
rect 48463 19594 48849 19613
rect 63583 19699 63969 19718
rect 63583 19676 63649 19699
rect 63735 19676 63817 19699
rect 63903 19676 63969 19699
rect 63583 19636 63592 19676
rect 63632 19636 63649 19676
rect 63735 19636 63756 19676
rect 63796 19636 63817 19676
rect 63903 19636 63920 19676
rect 63960 19636 63969 19676
rect 63583 19613 63649 19636
rect 63735 19613 63817 19636
rect 63903 19613 63969 19636
rect 63583 19594 63969 19613
rect 78703 19699 79089 19718
rect 78703 19676 78769 19699
rect 78855 19676 78937 19699
rect 79023 19676 79089 19699
rect 78703 19636 78712 19676
rect 78752 19636 78769 19676
rect 78855 19636 78876 19676
rect 78916 19636 78937 19676
rect 79023 19636 79040 19676
rect 79080 19636 79089 19676
rect 78703 19613 78769 19636
rect 78855 19613 78937 19636
rect 79023 19613 79089 19636
rect 78703 19594 79089 19613
rect 93823 19699 94209 19718
rect 93823 19676 93889 19699
rect 93975 19676 94057 19699
rect 94143 19676 94209 19699
rect 93823 19636 93832 19676
rect 93872 19636 93889 19676
rect 93975 19636 93996 19676
rect 94036 19636 94057 19676
rect 94143 19636 94160 19676
rect 94200 19636 94209 19676
rect 93823 19613 93889 19636
rect 93975 19613 94057 19636
rect 94143 19613 94209 19636
rect 93823 19594 94209 19613
rect 4343 18943 4729 18962
rect 4343 18920 4409 18943
rect 4495 18920 4577 18943
rect 4663 18920 4729 18943
rect 4343 18880 4352 18920
rect 4392 18880 4409 18920
rect 4495 18880 4516 18920
rect 4556 18880 4577 18920
rect 4663 18880 4680 18920
rect 4720 18880 4729 18920
rect 4343 18857 4409 18880
rect 4495 18857 4577 18880
rect 4663 18857 4729 18880
rect 4343 18838 4729 18857
rect 19463 18943 19849 18962
rect 19463 18920 19529 18943
rect 19615 18920 19697 18943
rect 19783 18920 19849 18943
rect 19463 18880 19472 18920
rect 19512 18880 19529 18920
rect 19615 18880 19636 18920
rect 19676 18880 19697 18920
rect 19783 18880 19800 18920
rect 19840 18880 19849 18920
rect 19463 18857 19529 18880
rect 19615 18857 19697 18880
rect 19783 18857 19849 18880
rect 19463 18838 19849 18857
rect 34583 18943 34969 18962
rect 34583 18920 34649 18943
rect 34735 18920 34817 18943
rect 34903 18920 34969 18943
rect 34583 18880 34592 18920
rect 34632 18880 34649 18920
rect 34735 18880 34756 18920
rect 34796 18880 34817 18920
rect 34903 18880 34920 18920
rect 34960 18880 34969 18920
rect 34583 18857 34649 18880
rect 34735 18857 34817 18880
rect 34903 18857 34969 18880
rect 34583 18838 34969 18857
rect 49703 18943 50089 18962
rect 49703 18920 49769 18943
rect 49855 18920 49937 18943
rect 50023 18920 50089 18943
rect 49703 18880 49712 18920
rect 49752 18880 49769 18920
rect 49855 18880 49876 18920
rect 49916 18880 49937 18920
rect 50023 18880 50040 18920
rect 50080 18880 50089 18920
rect 49703 18857 49769 18880
rect 49855 18857 49937 18880
rect 50023 18857 50089 18880
rect 49703 18838 50089 18857
rect 64823 18943 65209 18962
rect 64823 18920 64889 18943
rect 64975 18920 65057 18943
rect 65143 18920 65209 18943
rect 64823 18880 64832 18920
rect 64872 18880 64889 18920
rect 64975 18880 64996 18920
rect 65036 18880 65057 18920
rect 65143 18880 65160 18920
rect 65200 18880 65209 18920
rect 64823 18857 64889 18880
rect 64975 18857 65057 18880
rect 65143 18857 65209 18880
rect 64823 18838 65209 18857
rect 79943 18943 80329 18962
rect 79943 18920 80009 18943
rect 80095 18920 80177 18943
rect 80263 18920 80329 18943
rect 79943 18880 79952 18920
rect 79992 18880 80009 18920
rect 80095 18880 80116 18920
rect 80156 18880 80177 18920
rect 80263 18880 80280 18920
rect 80320 18880 80329 18920
rect 79943 18857 80009 18880
rect 80095 18857 80177 18880
rect 80263 18857 80329 18880
rect 79943 18838 80329 18857
rect 95063 18943 95449 18962
rect 95063 18920 95129 18943
rect 95215 18920 95297 18943
rect 95383 18920 95449 18943
rect 95063 18880 95072 18920
rect 95112 18880 95129 18920
rect 95215 18880 95236 18920
rect 95276 18880 95297 18920
rect 95383 18880 95400 18920
rect 95440 18880 95449 18920
rect 95063 18857 95129 18880
rect 95215 18857 95297 18880
rect 95383 18857 95449 18880
rect 95063 18838 95449 18857
rect 3103 18187 3489 18206
rect 3103 18164 3169 18187
rect 3255 18164 3337 18187
rect 3423 18164 3489 18187
rect 3103 18124 3112 18164
rect 3152 18124 3169 18164
rect 3255 18124 3276 18164
rect 3316 18124 3337 18164
rect 3423 18124 3440 18164
rect 3480 18124 3489 18164
rect 3103 18101 3169 18124
rect 3255 18101 3337 18124
rect 3423 18101 3489 18124
rect 3103 18082 3489 18101
rect 18223 18187 18609 18206
rect 18223 18164 18289 18187
rect 18375 18164 18457 18187
rect 18543 18164 18609 18187
rect 18223 18124 18232 18164
rect 18272 18124 18289 18164
rect 18375 18124 18396 18164
rect 18436 18124 18457 18164
rect 18543 18124 18560 18164
rect 18600 18124 18609 18164
rect 18223 18101 18289 18124
rect 18375 18101 18457 18124
rect 18543 18101 18609 18124
rect 18223 18082 18609 18101
rect 33343 18187 33729 18206
rect 33343 18164 33409 18187
rect 33495 18164 33577 18187
rect 33663 18164 33729 18187
rect 33343 18124 33352 18164
rect 33392 18124 33409 18164
rect 33495 18124 33516 18164
rect 33556 18124 33577 18164
rect 33663 18124 33680 18164
rect 33720 18124 33729 18164
rect 33343 18101 33409 18124
rect 33495 18101 33577 18124
rect 33663 18101 33729 18124
rect 33343 18082 33729 18101
rect 48463 18187 48849 18206
rect 48463 18164 48529 18187
rect 48615 18164 48697 18187
rect 48783 18164 48849 18187
rect 48463 18124 48472 18164
rect 48512 18124 48529 18164
rect 48615 18124 48636 18164
rect 48676 18124 48697 18164
rect 48783 18124 48800 18164
rect 48840 18124 48849 18164
rect 48463 18101 48529 18124
rect 48615 18101 48697 18124
rect 48783 18101 48849 18124
rect 48463 18082 48849 18101
rect 63583 18187 63969 18206
rect 63583 18164 63649 18187
rect 63735 18164 63817 18187
rect 63903 18164 63969 18187
rect 63583 18124 63592 18164
rect 63632 18124 63649 18164
rect 63735 18124 63756 18164
rect 63796 18124 63817 18164
rect 63903 18124 63920 18164
rect 63960 18124 63969 18164
rect 63583 18101 63649 18124
rect 63735 18101 63817 18124
rect 63903 18101 63969 18124
rect 63583 18082 63969 18101
rect 78703 18187 79089 18206
rect 78703 18164 78769 18187
rect 78855 18164 78937 18187
rect 79023 18164 79089 18187
rect 78703 18124 78712 18164
rect 78752 18124 78769 18164
rect 78855 18124 78876 18164
rect 78916 18124 78937 18164
rect 79023 18124 79040 18164
rect 79080 18124 79089 18164
rect 78703 18101 78769 18124
rect 78855 18101 78937 18124
rect 79023 18101 79089 18124
rect 78703 18082 79089 18101
rect 93823 18187 94209 18206
rect 93823 18164 93889 18187
rect 93975 18164 94057 18187
rect 94143 18164 94209 18187
rect 93823 18124 93832 18164
rect 93872 18124 93889 18164
rect 93975 18124 93996 18164
rect 94036 18124 94057 18164
rect 94143 18124 94160 18164
rect 94200 18124 94209 18164
rect 93823 18101 93889 18124
rect 93975 18101 94057 18124
rect 94143 18101 94209 18124
rect 93823 18082 94209 18101
rect 4343 17431 4729 17450
rect 4343 17408 4409 17431
rect 4495 17408 4577 17431
rect 4663 17408 4729 17431
rect 4343 17368 4352 17408
rect 4392 17368 4409 17408
rect 4495 17368 4516 17408
rect 4556 17368 4577 17408
rect 4663 17368 4680 17408
rect 4720 17368 4729 17408
rect 4343 17345 4409 17368
rect 4495 17345 4577 17368
rect 4663 17345 4729 17368
rect 4343 17326 4729 17345
rect 19463 17431 19849 17450
rect 19463 17408 19529 17431
rect 19615 17408 19697 17431
rect 19783 17408 19849 17431
rect 19463 17368 19472 17408
rect 19512 17368 19529 17408
rect 19615 17368 19636 17408
rect 19676 17368 19697 17408
rect 19783 17368 19800 17408
rect 19840 17368 19849 17408
rect 19463 17345 19529 17368
rect 19615 17345 19697 17368
rect 19783 17345 19849 17368
rect 19463 17326 19849 17345
rect 34583 17431 34969 17450
rect 34583 17408 34649 17431
rect 34735 17408 34817 17431
rect 34903 17408 34969 17431
rect 34583 17368 34592 17408
rect 34632 17368 34649 17408
rect 34735 17368 34756 17408
rect 34796 17368 34817 17408
rect 34903 17368 34920 17408
rect 34960 17368 34969 17408
rect 34583 17345 34649 17368
rect 34735 17345 34817 17368
rect 34903 17345 34969 17368
rect 34583 17326 34969 17345
rect 49703 17431 50089 17450
rect 49703 17408 49769 17431
rect 49855 17408 49937 17431
rect 50023 17408 50089 17431
rect 49703 17368 49712 17408
rect 49752 17368 49769 17408
rect 49855 17368 49876 17408
rect 49916 17368 49937 17408
rect 50023 17368 50040 17408
rect 50080 17368 50089 17408
rect 49703 17345 49769 17368
rect 49855 17345 49937 17368
rect 50023 17345 50089 17368
rect 49703 17326 50089 17345
rect 64823 17431 65209 17450
rect 64823 17408 64889 17431
rect 64975 17408 65057 17431
rect 65143 17408 65209 17431
rect 64823 17368 64832 17408
rect 64872 17368 64889 17408
rect 64975 17368 64996 17408
rect 65036 17368 65057 17408
rect 65143 17368 65160 17408
rect 65200 17368 65209 17408
rect 64823 17345 64889 17368
rect 64975 17345 65057 17368
rect 65143 17345 65209 17368
rect 64823 17326 65209 17345
rect 79943 17431 80329 17450
rect 79943 17408 80009 17431
rect 80095 17408 80177 17431
rect 80263 17408 80329 17431
rect 79943 17368 79952 17408
rect 79992 17368 80009 17408
rect 80095 17368 80116 17408
rect 80156 17368 80177 17408
rect 80263 17368 80280 17408
rect 80320 17368 80329 17408
rect 79943 17345 80009 17368
rect 80095 17345 80177 17368
rect 80263 17345 80329 17368
rect 79943 17326 80329 17345
rect 95063 17431 95449 17450
rect 95063 17408 95129 17431
rect 95215 17408 95297 17431
rect 95383 17408 95449 17431
rect 95063 17368 95072 17408
rect 95112 17368 95129 17408
rect 95215 17368 95236 17408
rect 95276 17368 95297 17408
rect 95383 17368 95400 17408
rect 95440 17368 95449 17408
rect 95063 17345 95129 17368
rect 95215 17345 95297 17368
rect 95383 17345 95449 17368
rect 95063 17326 95449 17345
rect 3103 16675 3489 16694
rect 3103 16652 3169 16675
rect 3255 16652 3337 16675
rect 3423 16652 3489 16675
rect 3103 16612 3112 16652
rect 3152 16612 3169 16652
rect 3255 16612 3276 16652
rect 3316 16612 3337 16652
rect 3423 16612 3440 16652
rect 3480 16612 3489 16652
rect 3103 16589 3169 16612
rect 3255 16589 3337 16612
rect 3423 16589 3489 16612
rect 3103 16570 3489 16589
rect 18223 16675 18609 16694
rect 18223 16652 18289 16675
rect 18375 16652 18457 16675
rect 18543 16652 18609 16675
rect 18223 16612 18232 16652
rect 18272 16612 18289 16652
rect 18375 16612 18396 16652
rect 18436 16612 18457 16652
rect 18543 16612 18560 16652
rect 18600 16612 18609 16652
rect 18223 16589 18289 16612
rect 18375 16589 18457 16612
rect 18543 16589 18609 16612
rect 18223 16570 18609 16589
rect 33343 16675 33729 16694
rect 33343 16652 33409 16675
rect 33495 16652 33577 16675
rect 33663 16652 33729 16675
rect 33343 16612 33352 16652
rect 33392 16612 33409 16652
rect 33495 16612 33516 16652
rect 33556 16612 33577 16652
rect 33663 16612 33680 16652
rect 33720 16612 33729 16652
rect 33343 16589 33409 16612
rect 33495 16589 33577 16612
rect 33663 16589 33729 16612
rect 33343 16570 33729 16589
rect 48463 16675 48849 16694
rect 48463 16652 48529 16675
rect 48615 16652 48697 16675
rect 48783 16652 48849 16675
rect 48463 16612 48472 16652
rect 48512 16612 48529 16652
rect 48615 16612 48636 16652
rect 48676 16612 48697 16652
rect 48783 16612 48800 16652
rect 48840 16612 48849 16652
rect 48463 16589 48529 16612
rect 48615 16589 48697 16612
rect 48783 16589 48849 16612
rect 48463 16570 48849 16589
rect 63583 16675 63969 16694
rect 63583 16652 63649 16675
rect 63735 16652 63817 16675
rect 63903 16652 63969 16675
rect 63583 16612 63592 16652
rect 63632 16612 63649 16652
rect 63735 16612 63756 16652
rect 63796 16612 63817 16652
rect 63903 16612 63920 16652
rect 63960 16612 63969 16652
rect 63583 16589 63649 16612
rect 63735 16589 63817 16612
rect 63903 16589 63969 16612
rect 63583 16570 63969 16589
rect 78703 16675 79089 16694
rect 78703 16652 78769 16675
rect 78855 16652 78937 16675
rect 79023 16652 79089 16675
rect 78703 16612 78712 16652
rect 78752 16612 78769 16652
rect 78855 16612 78876 16652
rect 78916 16612 78937 16652
rect 79023 16612 79040 16652
rect 79080 16612 79089 16652
rect 78703 16589 78769 16612
rect 78855 16589 78937 16612
rect 79023 16589 79089 16612
rect 78703 16570 79089 16589
rect 93823 16675 94209 16694
rect 93823 16652 93889 16675
rect 93975 16652 94057 16675
rect 94143 16652 94209 16675
rect 93823 16612 93832 16652
rect 93872 16612 93889 16652
rect 93975 16612 93996 16652
rect 94036 16612 94057 16652
rect 94143 16612 94160 16652
rect 94200 16612 94209 16652
rect 93823 16589 93889 16612
rect 93975 16589 94057 16612
rect 94143 16589 94209 16612
rect 93823 16570 94209 16589
rect 4343 15919 4729 15938
rect 4343 15896 4409 15919
rect 4495 15896 4577 15919
rect 4663 15896 4729 15919
rect 4343 15856 4352 15896
rect 4392 15856 4409 15896
rect 4495 15856 4516 15896
rect 4556 15856 4577 15896
rect 4663 15856 4680 15896
rect 4720 15856 4729 15896
rect 4343 15833 4409 15856
rect 4495 15833 4577 15856
rect 4663 15833 4729 15856
rect 4343 15814 4729 15833
rect 19463 15919 19849 15938
rect 19463 15896 19529 15919
rect 19615 15896 19697 15919
rect 19783 15896 19849 15919
rect 19463 15856 19472 15896
rect 19512 15856 19529 15896
rect 19615 15856 19636 15896
rect 19676 15856 19697 15896
rect 19783 15856 19800 15896
rect 19840 15856 19849 15896
rect 19463 15833 19529 15856
rect 19615 15833 19697 15856
rect 19783 15833 19849 15856
rect 19463 15814 19849 15833
rect 34583 15919 34969 15938
rect 34583 15896 34649 15919
rect 34735 15896 34817 15919
rect 34903 15896 34969 15919
rect 34583 15856 34592 15896
rect 34632 15856 34649 15896
rect 34735 15856 34756 15896
rect 34796 15856 34817 15896
rect 34903 15856 34920 15896
rect 34960 15856 34969 15896
rect 34583 15833 34649 15856
rect 34735 15833 34817 15856
rect 34903 15833 34969 15856
rect 34583 15814 34969 15833
rect 49703 15919 50089 15938
rect 49703 15896 49769 15919
rect 49855 15896 49937 15919
rect 50023 15896 50089 15919
rect 49703 15856 49712 15896
rect 49752 15856 49769 15896
rect 49855 15856 49876 15896
rect 49916 15856 49937 15896
rect 50023 15856 50040 15896
rect 50080 15856 50089 15896
rect 49703 15833 49769 15856
rect 49855 15833 49937 15856
rect 50023 15833 50089 15856
rect 49703 15814 50089 15833
rect 64823 15919 65209 15938
rect 64823 15896 64889 15919
rect 64975 15896 65057 15919
rect 65143 15896 65209 15919
rect 64823 15856 64832 15896
rect 64872 15856 64889 15896
rect 64975 15856 64996 15896
rect 65036 15856 65057 15896
rect 65143 15856 65160 15896
rect 65200 15856 65209 15896
rect 64823 15833 64889 15856
rect 64975 15833 65057 15856
rect 65143 15833 65209 15856
rect 64823 15814 65209 15833
rect 79943 15919 80329 15938
rect 79943 15896 80009 15919
rect 80095 15896 80177 15919
rect 80263 15896 80329 15919
rect 79943 15856 79952 15896
rect 79992 15856 80009 15896
rect 80095 15856 80116 15896
rect 80156 15856 80177 15896
rect 80263 15856 80280 15896
rect 80320 15856 80329 15896
rect 79943 15833 80009 15856
rect 80095 15833 80177 15856
rect 80263 15833 80329 15856
rect 79943 15814 80329 15833
rect 95063 15919 95449 15938
rect 95063 15896 95129 15919
rect 95215 15896 95297 15919
rect 95383 15896 95449 15919
rect 95063 15856 95072 15896
rect 95112 15856 95129 15896
rect 95215 15856 95236 15896
rect 95276 15856 95297 15896
rect 95383 15856 95400 15896
rect 95440 15856 95449 15896
rect 95063 15833 95129 15856
rect 95215 15833 95297 15856
rect 95383 15833 95449 15856
rect 95063 15814 95449 15833
rect 3103 15163 3489 15182
rect 3103 15140 3169 15163
rect 3255 15140 3337 15163
rect 3423 15140 3489 15163
rect 3103 15100 3112 15140
rect 3152 15100 3169 15140
rect 3255 15100 3276 15140
rect 3316 15100 3337 15140
rect 3423 15100 3440 15140
rect 3480 15100 3489 15140
rect 3103 15077 3169 15100
rect 3255 15077 3337 15100
rect 3423 15077 3489 15100
rect 3103 15058 3489 15077
rect 18223 15163 18609 15182
rect 18223 15140 18289 15163
rect 18375 15140 18457 15163
rect 18543 15140 18609 15163
rect 18223 15100 18232 15140
rect 18272 15100 18289 15140
rect 18375 15100 18396 15140
rect 18436 15100 18457 15140
rect 18543 15100 18560 15140
rect 18600 15100 18609 15140
rect 18223 15077 18289 15100
rect 18375 15077 18457 15100
rect 18543 15077 18609 15100
rect 18223 15058 18609 15077
rect 33343 15163 33729 15182
rect 33343 15140 33409 15163
rect 33495 15140 33577 15163
rect 33663 15140 33729 15163
rect 33343 15100 33352 15140
rect 33392 15100 33409 15140
rect 33495 15100 33516 15140
rect 33556 15100 33577 15140
rect 33663 15100 33680 15140
rect 33720 15100 33729 15140
rect 33343 15077 33409 15100
rect 33495 15077 33577 15100
rect 33663 15077 33729 15100
rect 33343 15058 33729 15077
rect 48463 15163 48849 15182
rect 48463 15140 48529 15163
rect 48615 15140 48697 15163
rect 48783 15140 48849 15163
rect 48463 15100 48472 15140
rect 48512 15100 48529 15140
rect 48615 15100 48636 15140
rect 48676 15100 48697 15140
rect 48783 15100 48800 15140
rect 48840 15100 48849 15140
rect 48463 15077 48529 15100
rect 48615 15077 48697 15100
rect 48783 15077 48849 15100
rect 48463 15058 48849 15077
rect 63583 15163 63969 15182
rect 63583 15140 63649 15163
rect 63735 15140 63817 15163
rect 63903 15140 63969 15163
rect 63583 15100 63592 15140
rect 63632 15100 63649 15140
rect 63735 15100 63756 15140
rect 63796 15100 63817 15140
rect 63903 15100 63920 15140
rect 63960 15100 63969 15140
rect 63583 15077 63649 15100
rect 63735 15077 63817 15100
rect 63903 15077 63969 15100
rect 63583 15058 63969 15077
rect 78703 15163 79089 15182
rect 78703 15140 78769 15163
rect 78855 15140 78937 15163
rect 79023 15140 79089 15163
rect 78703 15100 78712 15140
rect 78752 15100 78769 15140
rect 78855 15100 78876 15140
rect 78916 15100 78937 15140
rect 79023 15100 79040 15140
rect 79080 15100 79089 15140
rect 78703 15077 78769 15100
rect 78855 15077 78937 15100
rect 79023 15077 79089 15100
rect 78703 15058 79089 15077
rect 93823 15163 94209 15182
rect 93823 15140 93889 15163
rect 93975 15140 94057 15163
rect 94143 15140 94209 15163
rect 93823 15100 93832 15140
rect 93872 15100 93889 15140
rect 93975 15100 93996 15140
rect 94036 15100 94057 15140
rect 94143 15100 94160 15140
rect 94200 15100 94209 15140
rect 93823 15077 93889 15100
rect 93975 15077 94057 15100
rect 94143 15077 94209 15100
rect 93823 15058 94209 15077
rect 4343 14407 4729 14426
rect 4343 14384 4409 14407
rect 4495 14384 4577 14407
rect 4663 14384 4729 14407
rect 4343 14344 4352 14384
rect 4392 14344 4409 14384
rect 4495 14344 4516 14384
rect 4556 14344 4577 14384
rect 4663 14344 4680 14384
rect 4720 14344 4729 14384
rect 4343 14321 4409 14344
rect 4495 14321 4577 14344
rect 4663 14321 4729 14344
rect 4343 14302 4729 14321
rect 19463 14407 19849 14426
rect 19463 14384 19529 14407
rect 19615 14384 19697 14407
rect 19783 14384 19849 14407
rect 19463 14344 19472 14384
rect 19512 14344 19529 14384
rect 19615 14344 19636 14384
rect 19676 14344 19697 14384
rect 19783 14344 19800 14384
rect 19840 14344 19849 14384
rect 19463 14321 19529 14344
rect 19615 14321 19697 14344
rect 19783 14321 19849 14344
rect 19463 14302 19849 14321
rect 34583 14407 34969 14426
rect 34583 14384 34649 14407
rect 34735 14384 34817 14407
rect 34903 14384 34969 14407
rect 34583 14344 34592 14384
rect 34632 14344 34649 14384
rect 34735 14344 34756 14384
rect 34796 14344 34817 14384
rect 34903 14344 34920 14384
rect 34960 14344 34969 14384
rect 34583 14321 34649 14344
rect 34735 14321 34817 14344
rect 34903 14321 34969 14344
rect 34583 14302 34969 14321
rect 49703 14407 50089 14426
rect 49703 14384 49769 14407
rect 49855 14384 49937 14407
rect 50023 14384 50089 14407
rect 49703 14344 49712 14384
rect 49752 14344 49769 14384
rect 49855 14344 49876 14384
rect 49916 14344 49937 14384
rect 50023 14344 50040 14384
rect 50080 14344 50089 14384
rect 49703 14321 49769 14344
rect 49855 14321 49937 14344
rect 50023 14321 50089 14344
rect 49703 14302 50089 14321
rect 64823 14407 65209 14426
rect 64823 14384 64889 14407
rect 64975 14384 65057 14407
rect 65143 14384 65209 14407
rect 64823 14344 64832 14384
rect 64872 14344 64889 14384
rect 64975 14344 64996 14384
rect 65036 14344 65057 14384
rect 65143 14344 65160 14384
rect 65200 14344 65209 14384
rect 64823 14321 64889 14344
rect 64975 14321 65057 14344
rect 65143 14321 65209 14344
rect 64823 14302 65209 14321
rect 79943 14407 80329 14426
rect 79943 14384 80009 14407
rect 80095 14384 80177 14407
rect 80263 14384 80329 14407
rect 79943 14344 79952 14384
rect 79992 14344 80009 14384
rect 80095 14344 80116 14384
rect 80156 14344 80177 14384
rect 80263 14344 80280 14384
rect 80320 14344 80329 14384
rect 79943 14321 80009 14344
rect 80095 14321 80177 14344
rect 80263 14321 80329 14344
rect 79943 14302 80329 14321
rect 95063 14407 95449 14426
rect 95063 14384 95129 14407
rect 95215 14384 95297 14407
rect 95383 14384 95449 14407
rect 95063 14344 95072 14384
rect 95112 14344 95129 14384
rect 95215 14344 95236 14384
rect 95276 14344 95297 14384
rect 95383 14344 95400 14384
rect 95440 14344 95449 14384
rect 95063 14321 95129 14344
rect 95215 14321 95297 14344
rect 95383 14321 95449 14344
rect 95063 14302 95449 14321
rect 3103 13651 3489 13670
rect 3103 13628 3169 13651
rect 3255 13628 3337 13651
rect 3423 13628 3489 13651
rect 3103 13588 3112 13628
rect 3152 13588 3169 13628
rect 3255 13588 3276 13628
rect 3316 13588 3337 13628
rect 3423 13588 3440 13628
rect 3480 13588 3489 13628
rect 3103 13565 3169 13588
rect 3255 13565 3337 13588
rect 3423 13565 3489 13588
rect 3103 13546 3489 13565
rect 18223 13651 18609 13670
rect 18223 13628 18289 13651
rect 18375 13628 18457 13651
rect 18543 13628 18609 13651
rect 18223 13588 18232 13628
rect 18272 13588 18289 13628
rect 18375 13588 18396 13628
rect 18436 13588 18457 13628
rect 18543 13588 18560 13628
rect 18600 13588 18609 13628
rect 18223 13565 18289 13588
rect 18375 13565 18457 13588
rect 18543 13565 18609 13588
rect 18223 13546 18609 13565
rect 33343 13651 33729 13670
rect 33343 13628 33409 13651
rect 33495 13628 33577 13651
rect 33663 13628 33729 13651
rect 33343 13588 33352 13628
rect 33392 13588 33409 13628
rect 33495 13588 33516 13628
rect 33556 13588 33577 13628
rect 33663 13588 33680 13628
rect 33720 13588 33729 13628
rect 33343 13565 33409 13588
rect 33495 13565 33577 13588
rect 33663 13565 33729 13588
rect 33343 13546 33729 13565
rect 48463 13651 48849 13670
rect 48463 13628 48529 13651
rect 48615 13628 48697 13651
rect 48783 13628 48849 13651
rect 48463 13588 48472 13628
rect 48512 13588 48529 13628
rect 48615 13588 48636 13628
rect 48676 13588 48697 13628
rect 48783 13588 48800 13628
rect 48840 13588 48849 13628
rect 48463 13565 48529 13588
rect 48615 13565 48697 13588
rect 48783 13565 48849 13588
rect 48463 13546 48849 13565
rect 63583 13651 63969 13670
rect 63583 13628 63649 13651
rect 63735 13628 63817 13651
rect 63903 13628 63969 13651
rect 63583 13588 63592 13628
rect 63632 13588 63649 13628
rect 63735 13588 63756 13628
rect 63796 13588 63817 13628
rect 63903 13588 63920 13628
rect 63960 13588 63969 13628
rect 63583 13565 63649 13588
rect 63735 13565 63817 13588
rect 63903 13565 63969 13588
rect 63583 13546 63969 13565
rect 78703 13651 79089 13670
rect 78703 13628 78769 13651
rect 78855 13628 78937 13651
rect 79023 13628 79089 13651
rect 78703 13588 78712 13628
rect 78752 13588 78769 13628
rect 78855 13588 78876 13628
rect 78916 13588 78937 13628
rect 79023 13588 79040 13628
rect 79080 13588 79089 13628
rect 78703 13565 78769 13588
rect 78855 13565 78937 13588
rect 79023 13565 79089 13588
rect 78703 13546 79089 13565
rect 93823 13651 94209 13670
rect 93823 13628 93889 13651
rect 93975 13628 94057 13651
rect 94143 13628 94209 13651
rect 93823 13588 93832 13628
rect 93872 13588 93889 13628
rect 93975 13588 93996 13628
rect 94036 13588 94057 13628
rect 94143 13588 94160 13628
rect 94200 13588 94209 13628
rect 93823 13565 93889 13588
rect 93975 13565 94057 13588
rect 94143 13565 94209 13588
rect 93823 13546 94209 13565
rect 4343 12895 4729 12914
rect 4343 12872 4409 12895
rect 4495 12872 4577 12895
rect 4663 12872 4729 12895
rect 4343 12832 4352 12872
rect 4392 12832 4409 12872
rect 4495 12832 4516 12872
rect 4556 12832 4577 12872
rect 4663 12832 4680 12872
rect 4720 12832 4729 12872
rect 4343 12809 4409 12832
rect 4495 12809 4577 12832
rect 4663 12809 4729 12832
rect 4343 12790 4729 12809
rect 19463 12895 19849 12914
rect 19463 12872 19529 12895
rect 19615 12872 19697 12895
rect 19783 12872 19849 12895
rect 19463 12832 19472 12872
rect 19512 12832 19529 12872
rect 19615 12832 19636 12872
rect 19676 12832 19697 12872
rect 19783 12832 19800 12872
rect 19840 12832 19849 12872
rect 19463 12809 19529 12832
rect 19615 12809 19697 12832
rect 19783 12809 19849 12832
rect 19463 12790 19849 12809
rect 34583 12895 34969 12914
rect 34583 12872 34649 12895
rect 34735 12872 34817 12895
rect 34903 12872 34969 12895
rect 34583 12832 34592 12872
rect 34632 12832 34649 12872
rect 34735 12832 34756 12872
rect 34796 12832 34817 12872
rect 34903 12832 34920 12872
rect 34960 12832 34969 12872
rect 34583 12809 34649 12832
rect 34735 12809 34817 12832
rect 34903 12809 34969 12832
rect 34583 12790 34969 12809
rect 49703 12895 50089 12914
rect 49703 12872 49769 12895
rect 49855 12872 49937 12895
rect 50023 12872 50089 12895
rect 49703 12832 49712 12872
rect 49752 12832 49769 12872
rect 49855 12832 49876 12872
rect 49916 12832 49937 12872
rect 50023 12832 50040 12872
rect 50080 12832 50089 12872
rect 49703 12809 49769 12832
rect 49855 12809 49937 12832
rect 50023 12809 50089 12832
rect 49703 12790 50089 12809
rect 64823 12895 65209 12914
rect 64823 12872 64889 12895
rect 64975 12872 65057 12895
rect 65143 12872 65209 12895
rect 64823 12832 64832 12872
rect 64872 12832 64889 12872
rect 64975 12832 64996 12872
rect 65036 12832 65057 12872
rect 65143 12832 65160 12872
rect 65200 12832 65209 12872
rect 64823 12809 64889 12832
rect 64975 12809 65057 12832
rect 65143 12809 65209 12832
rect 64823 12790 65209 12809
rect 79943 12895 80329 12914
rect 79943 12872 80009 12895
rect 80095 12872 80177 12895
rect 80263 12872 80329 12895
rect 79943 12832 79952 12872
rect 79992 12832 80009 12872
rect 80095 12832 80116 12872
rect 80156 12832 80177 12872
rect 80263 12832 80280 12872
rect 80320 12832 80329 12872
rect 79943 12809 80009 12832
rect 80095 12809 80177 12832
rect 80263 12809 80329 12832
rect 79943 12790 80329 12809
rect 95063 12895 95449 12914
rect 95063 12872 95129 12895
rect 95215 12872 95297 12895
rect 95383 12872 95449 12895
rect 95063 12832 95072 12872
rect 95112 12832 95129 12872
rect 95215 12832 95236 12872
rect 95276 12832 95297 12872
rect 95383 12832 95400 12872
rect 95440 12832 95449 12872
rect 95063 12809 95129 12832
rect 95215 12809 95297 12832
rect 95383 12809 95449 12832
rect 95063 12790 95449 12809
rect 3103 12139 3489 12158
rect 3103 12116 3169 12139
rect 3255 12116 3337 12139
rect 3423 12116 3489 12139
rect 3103 12076 3112 12116
rect 3152 12076 3169 12116
rect 3255 12076 3276 12116
rect 3316 12076 3337 12116
rect 3423 12076 3440 12116
rect 3480 12076 3489 12116
rect 3103 12053 3169 12076
rect 3255 12053 3337 12076
rect 3423 12053 3489 12076
rect 3103 12034 3489 12053
rect 18223 12139 18609 12158
rect 18223 12116 18289 12139
rect 18375 12116 18457 12139
rect 18543 12116 18609 12139
rect 18223 12076 18232 12116
rect 18272 12076 18289 12116
rect 18375 12076 18396 12116
rect 18436 12076 18457 12116
rect 18543 12076 18560 12116
rect 18600 12076 18609 12116
rect 18223 12053 18289 12076
rect 18375 12053 18457 12076
rect 18543 12053 18609 12076
rect 18223 12034 18609 12053
rect 33343 12139 33729 12158
rect 33343 12116 33409 12139
rect 33495 12116 33577 12139
rect 33663 12116 33729 12139
rect 33343 12076 33352 12116
rect 33392 12076 33409 12116
rect 33495 12076 33516 12116
rect 33556 12076 33577 12116
rect 33663 12076 33680 12116
rect 33720 12076 33729 12116
rect 33343 12053 33409 12076
rect 33495 12053 33577 12076
rect 33663 12053 33729 12076
rect 33343 12034 33729 12053
rect 48463 12139 48849 12158
rect 48463 12116 48529 12139
rect 48615 12116 48697 12139
rect 48783 12116 48849 12139
rect 48463 12076 48472 12116
rect 48512 12076 48529 12116
rect 48615 12076 48636 12116
rect 48676 12076 48697 12116
rect 48783 12076 48800 12116
rect 48840 12076 48849 12116
rect 48463 12053 48529 12076
rect 48615 12053 48697 12076
rect 48783 12053 48849 12076
rect 48463 12034 48849 12053
rect 63583 12139 63969 12158
rect 63583 12116 63649 12139
rect 63735 12116 63817 12139
rect 63903 12116 63969 12139
rect 63583 12076 63592 12116
rect 63632 12076 63649 12116
rect 63735 12076 63756 12116
rect 63796 12076 63817 12116
rect 63903 12076 63920 12116
rect 63960 12076 63969 12116
rect 63583 12053 63649 12076
rect 63735 12053 63817 12076
rect 63903 12053 63969 12076
rect 63583 12034 63969 12053
rect 78703 12139 79089 12158
rect 78703 12116 78769 12139
rect 78855 12116 78937 12139
rect 79023 12116 79089 12139
rect 78703 12076 78712 12116
rect 78752 12076 78769 12116
rect 78855 12076 78876 12116
rect 78916 12076 78937 12116
rect 79023 12076 79040 12116
rect 79080 12076 79089 12116
rect 78703 12053 78769 12076
rect 78855 12053 78937 12076
rect 79023 12053 79089 12076
rect 78703 12034 79089 12053
rect 93823 12139 94209 12158
rect 93823 12116 93889 12139
rect 93975 12116 94057 12139
rect 94143 12116 94209 12139
rect 93823 12076 93832 12116
rect 93872 12076 93889 12116
rect 93975 12076 93996 12116
rect 94036 12076 94057 12116
rect 94143 12076 94160 12116
rect 94200 12076 94209 12116
rect 93823 12053 93889 12076
rect 93975 12053 94057 12076
rect 94143 12053 94209 12076
rect 93823 12034 94209 12053
rect 4343 11383 4729 11402
rect 4343 11360 4409 11383
rect 4495 11360 4577 11383
rect 4663 11360 4729 11383
rect 4343 11320 4352 11360
rect 4392 11320 4409 11360
rect 4495 11320 4516 11360
rect 4556 11320 4577 11360
rect 4663 11320 4680 11360
rect 4720 11320 4729 11360
rect 4343 11297 4409 11320
rect 4495 11297 4577 11320
rect 4663 11297 4729 11320
rect 4343 11278 4729 11297
rect 19463 11383 19849 11402
rect 19463 11360 19529 11383
rect 19615 11360 19697 11383
rect 19783 11360 19849 11383
rect 19463 11320 19472 11360
rect 19512 11320 19529 11360
rect 19615 11320 19636 11360
rect 19676 11320 19697 11360
rect 19783 11320 19800 11360
rect 19840 11320 19849 11360
rect 19463 11297 19529 11320
rect 19615 11297 19697 11320
rect 19783 11297 19849 11320
rect 19463 11278 19849 11297
rect 34583 11383 34969 11402
rect 34583 11360 34649 11383
rect 34735 11360 34817 11383
rect 34903 11360 34969 11383
rect 34583 11320 34592 11360
rect 34632 11320 34649 11360
rect 34735 11320 34756 11360
rect 34796 11320 34817 11360
rect 34903 11320 34920 11360
rect 34960 11320 34969 11360
rect 34583 11297 34649 11320
rect 34735 11297 34817 11320
rect 34903 11297 34969 11320
rect 34583 11278 34969 11297
rect 49703 11383 50089 11402
rect 49703 11360 49769 11383
rect 49855 11360 49937 11383
rect 50023 11360 50089 11383
rect 49703 11320 49712 11360
rect 49752 11320 49769 11360
rect 49855 11320 49876 11360
rect 49916 11320 49937 11360
rect 50023 11320 50040 11360
rect 50080 11320 50089 11360
rect 49703 11297 49769 11320
rect 49855 11297 49937 11320
rect 50023 11297 50089 11320
rect 49703 11278 50089 11297
rect 64823 11383 65209 11402
rect 64823 11360 64889 11383
rect 64975 11360 65057 11383
rect 65143 11360 65209 11383
rect 64823 11320 64832 11360
rect 64872 11320 64889 11360
rect 64975 11320 64996 11360
rect 65036 11320 65057 11360
rect 65143 11320 65160 11360
rect 65200 11320 65209 11360
rect 64823 11297 64889 11320
rect 64975 11297 65057 11320
rect 65143 11297 65209 11320
rect 64823 11278 65209 11297
rect 79943 11383 80329 11402
rect 79943 11360 80009 11383
rect 80095 11360 80177 11383
rect 80263 11360 80329 11383
rect 79943 11320 79952 11360
rect 79992 11320 80009 11360
rect 80095 11320 80116 11360
rect 80156 11320 80177 11360
rect 80263 11320 80280 11360
rect 80320 11320 80329 11360
rect 79943 11297 80009 11320
rect 80095 11297 80177 11320
rect 80263 11297 80329 11320
rect 79943 11278 80329 11297
rect 95063 11383 95449 11402
rect 95063 11360 95129 11383
rect 95215 11360 95297 11383
rect 95383 11360 95449 11383
rect 95063 11320 95072 11360
rect 95112 11320 95129 11360
rect 95215 11320 95236 11360
rect 95276 11320 95297 11360
rect 95383 11320 95400 11360
rect 95440 11320 95449 11360
rect 95063 11297 95129 11320
rect 95215 11297 95297 11320
rect 95383 11297 95449 11320
rect 95063 11278 95449 11297
rect 3103 10627 3489 10646
rect 3103 10604 3169 10627
rect 3255 10604 3337 10627
rect 3423 10604 3489 10627
rect 3103 10564 3112 10604
rect 3152 10564 3169 10604
rect 3255 10564 3276 10604
rect 3316 10564 3337 10604
rect 3423 10564 3440 10604
rect 3480 10564 3489 10604
rect 3103 10541 3169 10564
rect 3255 10541 3337 10564
rect 3423 10541 3489 10564
rect 3103 10522 3489 10541
rect 18223 10627 18609 10646
rect 18223 10604 18289 10627
rect 18375 10604 18457 10627
rect 18543 10604 18609 10627
rect 18223 10564 18232 10604
rect 18272 10564 18289 10604
rect 18375 10564 18396 10604
rect 18436 10564 18457 10604
rect 18543 10564 18560 10604
rect 18600 10564 18609 10604
rect 18223 10541 18289 10564
rect 18375 10541 18457 10564
rect 18543 10541 18609 10564
rect 18223 10522 18609 10541
rect 33343 10627 33729 10646
rect 33343 10604 33409 10627
rect 33495 10604 33577 10627
rect 33663 10604 33729 10627
rect 33343 10564 33352 10604
rect 33392 10564 33409 10604
rect 33495 10564 33516 10604
rect 33556 10564 33577 10604
rect 33663 10564 33680 10604
rect 33720 10564 33729 10604
rect 33343 10541 33409 10564
rect 33495 10541 33577 10564
rect 33663 10541 33729 10564
rect 33343 10522 33729 10541
rect 48463 10627 48849 10646
rect 48463 10604 48529 10627
rect 48615 10604 48697 10627
rect 48783 10604 48849 10627
rect 48463 10564 48472 10604
rect 48512 10564 48529 10604
rect 48615 10564 48636 10604
rect 48676 10564 48697 10604
rect 48783 10564 48800 10604
rect 48840 10564 48849 10604
rect 48463 10541 48529 10564
rect 48615 10541 48697 10564
rect 48783 10541 48849 10564
rect 48463 10522 48849 10541
rect 63583 10627 63969 10646
rect 63583 10604 63649 10627
rect 63735 10604 63817 10627
rect 63903 10604 63969 10627
rect 63583 10564 63592 10604
rect 63632 10564 63649 10604
rect 63735 10564 63756 10604
rect 63796 10564 63817 10604
rect 63903 10564 63920 10604
rect 63960 10564 63969 10604
rect 63583 10541 63649 10564
rect 63735 10541 63817 10564
rect 63903 10541 63969 10564
rect 63583 10522 63969 10541
rect 78703 10627 79089 10646
rect 78703 10604 78769 10627
rect 78855 10604 78937 10627
rect 79023 10604 79089 10627
rect 78703 10564 78712 10604
rect 78752 10564 78769 10604
rect 78855 10564 78876 10604
rect 78916 10564 78937 10604
rect 79023 10564 79040 10604
rect 79080 10564 79089 10604
rect 78703 10541 78769 10564
rect 78855 10541 78937 10564
rect 79023 10541 79089 10564
rect 78703 10522 79089 10541
rect 93823 10627 94209 10646
rect 93823 10604 93889 10627
rect 93975 10604 94057 10627
rect 94143 10604 94209 10627
rect 93823 10564 93832 10604
rect 93872 10564 93889 10604
rect 93975 10564 93996 10604
rect 94036 10564 94057 10604
rect 94143 10564 94160 10604
rect 94200 10564 94209 10604
rect 93823 10541 93889 10564
rect 93975 10541 94057 10564
rect 94143 10541 94209 10564
rect 93823 10522 94209 10541
rect 4343 9871 4729 9890
rect 4343 9848 4409 9871
rect 4495 9848 4577 9871
rect 4663 9848 4729 9871
rect 4343 9808 4352 9848
rect 4392 9808 4409 9848
rect 4495 9808 4516 9848
rect 4556 9808 4577 9848
rect 4663 9808 4680 9848
rect 4720 9808 4729 9848
rect 4343 9785 4409 9808
rect 4495 9785 4577 9808
rect 4663 9785 4729 9808
rect 4343 9766 4729 9785
rect 19463 9871 19849 9890
rect 19463 9848 19529 9871
rect 19615 9848 19697 9871
rect 19783 9848 19849 9871
rect 19463 9808 19472 9848
rect 19512 9808 19529 9848
rect 19615 9808 19636 9848
rect 19676 9808 19697 9848
rect 19783 9808 19800 9848
rect 19840 9808 19849 9848
rect 19463 9785 19529 9808
rect 19615 9785 19697 9808
rect 19783 9785 19849 9808
rect 19463 9766 19849 9785
rect 34583 9871 34969 9890
rect 34583 9848 34649 9871
rect 34735 9848 34817 9871
rect 34903 9848 34969 9871
rect 34583 9808 34592 9848
rect 34632 9808 34649 9848
rect 34735 9808 34756 9848
rect 34796 9808 34817 9848
rect 34903 9808 34920 9848
rect 34960 9808 34969 9848
rect 34583 9785 34649 9808
rect 34735 9785 34817 9808
rect 34903 9785 34969 9808
rect 34583 9766 34969 9785
rect 49703 9871 50089 9890
rect 49703 9848 49769 9871
rect 49855 9848 49937 9871
rect 50023 9848 50089 9871
rect 49703 9808 49712 9848
rect 49752 9808 49769 9848
rect 49855 9808 49876 9848
rect 49916 9808 49937 9848
rect 50023 9808 50040 9848
rect 50080 9808 50089 9848
rect 49703 9785 49769 9808
rect 49855 9785 49937 9808
rect 50023 9785 50089 9808
rect 49703 9766 50089 9785
rect 64823 9871 65209 9890
rect 64823 9848 64889 9871
rect 64975 9848 65057 9871
rect 65143 9848 65209 9871
rect 64823 9808 64832 9848
rect 64872 9808 64889 9848
rect 64975 9808 64996 9848
rect 65036 9808 65057 9848
rect 65143 9808 65160 9848
rect 65200 9808 65209 9848
rect 64823 9785 64889 9808
rect 64975 9785 65057 9808
rect 65143 9785 65209 9808
rect 64823 9766 65209 9785
rect 79943 9871 80329 9890
rect 79943 9848 80009 9871
rect 80095 9848 80177 9871
rect 80263 9848 80329 9871
rect 79943 9808 79952 9848
rect 79992 9808 80009 9848
rect 80095 9808 80116 9848
rect 80156 9808 80177 9848
rect 80263 9808 80280 9848
rect 80320 9808 80329 9848
rect 79943 9785 80009 9808
rect 80095 9785 80177 9808
rect 80263 9785 80329 9808
rect 79943 9766 80329 9785
rect 95063 9871 95449 9890
rect 95063 9848 95129 9871
rect 95215 9848 95297 9871
rect 95383 9848 95449 9871
rect 95063 9808 95072 9848
rect 95112 9808 95129 9848
rect 95215 9808 95236 9848
rect 95276 9808 95297 9848
rect 95383 9808 95400 9848
rect 95440 9808 95449 9848
rect 95063 9785 95129 9808
rect 95215 9785 95297 9808
rect 95383 9785 95449 9808
rect 95063 9766 95449 9785
rect 3103 9115 3489 9134
rect 3103 9092 3169 9115
rect 3255 9092 3337 9115
rect 3423 9092 3489 9115
rect 3103 9052 3112 9092
rect 3152 9052 3169 9092
rect 3255 9052 3276 9092
rect 3316 9052 3337 9092
rect 3423 9052 3440 9092
rect 3480 9052 3489 9092
rect 3103 9029 3169 9052
rect 3255 9029 3337 9052
rect 3423 9029 3489 9052
rect 3103 9010 3489 9029
rect 18223 9115 18609 9134
rect 18223 9092 18289 9115
rect 18375 9092 18457 9115
rect 18543 9092 18609 9115
rect 18223 9052 18232 9092
rect 18272 9052 18289 9092
rect 18375 9052 18396 9092
rect 18436 9052 18457 9092
rect 18543 9052 18560 9092
rect 18600 9052 18609 9092
rect 18223 9029 18289 9052
rect 18375 9029 18457 9052
rect 18543 9029 18609 9052
rect 18223 9010 18609 9029
rect 33343 9115 33729 9134
rect 33343 9092 33409 9115
rect 33495 9092 33577 9115
rect 33663 9092 33729 9115
rect 33343 9052 33352 9092
rect 33392 9052 33409 9092
rect 33495 9052 33516 9092
rect 33556 9052 33577 9092
rect 33663 9052 33680 9092
rect 33720 9052 33729 9092
rect 33343 9029 33409 9052
rect 33495 9029 33577 9052
rect 33663 9029 33729 9052
rect 33343 9010 33729 9029
rect 48463 9115 48849 9134
rect 48463 9092 48529 9115
rect 48615 9092 48697 9115
rect 48783 9092 48849 9115
rect 48463 9052 48472 9092
rect 48512 9052 48529 9092
rect 48615 9052 48636 9092
rect 48676 9052 48697 9092
rect 48783 9052 48800 9092
rect 48840 9052 48849 9092
rect 48463 9029 48529 9052
rect 48615 9029 48697 9052
rect 48783 9029 48849 9052
rect 48463 9010 48849 9029
rect 63583 9115 63969 9134
rect 63583 9092 63649 9115
rect 63735 9092 63817 9115
rect 63903 9092 63969 9115
rect 63583 9052 63592 9092
rect 63632 9052 63649 9092
rect 63735 9052 63756 9092
rect 63796 9052 63817 9092
rect 63903 9052 63920 9092
rect 63960 9052 63969 9092
rect 63583 9029 63649 9052
rect 63735 9029 63817 9052
rect 63903 9029 63969 9052
rect 63583 9010 63969 9029
rect 78703 9115 79089 9134
rect 78703 9092 78769 9115
rect 78855 9092 78937 9115
rect 79023 9092 79089 9115
rect 78703 9052 78712 9092
rect 78752 9052 78769 9092
rect 78855 9052 78876 9092
rect 78916 9052 78937 9092
rect 79023 9052 79040 9092
rect 79080 9052 79089 9092
rect 78703 9029 78769 9052
rect 78855 9029 78937 9052
rect 79023 9029 79089 9052
rect 78703 9010 79089 9029
rect 93823 9115 94209 9134
rect 93823 9092 93889 9115
rect 93975 9092 94057 9115
rect 94143 9092 94209 9115
rect 93823 9052 93832 9092
rect 93872 9052 93889 9092
rect 93975 9052 93996 9092
rect 94036 9052 94057 9092
rect 94143 9052 94160 9092
rect 94200 9052 94209 9092
rect 93823 9029 93889 9052
rect 93975 9029 94057 9052
rect 94143 9029 94209 9052
rect 93823 9010 94209 9029
rect 4343 8359 4729 8378
rect 4343 8336 4409 8359
rect 4495 8336 4577 8359
rect 4663 8336 4729 8359
rect 4343 8296 4352 8336
rect 4392 8296 4409 8336
rect 4495 8296 4516 8336
rect 4556 8296 4577 8336
rect 4663 8296 4680 8336
rect 4720 8296 4729 8336
rect 4343 8273 4409 8296
rect 4495 8273 4577 8296
rect 4663 8273 4729 8296
rect 4343 8254 4729 8273
rect 19463 8359 19849 8378
rect 19463 8336 19529 8359
rect 19615 8336 19697 8359
rect 19783 8336 19849 8359
rect 19463 8296 19472 8336
rect 19512 8296 19529 8336
rect 19615 8296 19636 8336
rect 19676 8296 19697 8336
rect 19783 8296 19800 8336
rect 19840 8296 19849 8336
rect 19463 8273 19529 8296
rect 19615 8273 19697 8296
rect 19783 8273 19849 8296
rect 19463 8254 19849 8273
rect 34583 8359 34969 8378
rect 34583 8336 34649 8359
rect 34735 8336 34817 8359
rect 34903 8336 34969 8359
rect 34583 8296 34592 8336
rect 34632 8296 34649 8336
rect 34735 8296 34756 8336
rect 34796 8296 34817 8336
rect 34903 8296 34920 8336
rect 34960 8296 34969 8336
rect 34583 8273 34649 8296
rect 34735 8273 34817 8296
rect 34903 8273 34969 8296
rect 34583 8254 34969 8273
rect 49703 8359 50089 8378
rect 49703 8336 49769 8359
rect 49855 8336 49937 8359
rect 50023 8336 50089 8359
rect 49703 8296 49712 8336
rect 49752 8296 49769 8336
rect 49855 8296 49876 8336
rect 49916 8296 49937 8336
rect 50023 8296 50040 8336
rect 50080 8296 50089 8336
rect 49703 8273 49769 8296
rect 49855 8273 49937 8296
rect 50023 8273 50089 8296
rect 49703 8254 50089 8273
rect 64823 8359 65209 8378
rect 64823 8336 64889 8359
rect 64975 8336 65057 8359
rect 65143 8336 65209 8359
rect 64823 8296 64832 8336
rect 64872 8296 64889 8336
rect 64975 8296 64996 8336
rect 65036 8296 65057 8336
rect 65143 8296 65160 8336
rect 65200 8296 65209 8336
rect 64823 8273 64889 8296
rect 64975 8273 65057 8296
rect 65143 8273 65209 8296
rect 64823 8254 65209 8273
rect 79943 8359 80329 8378
rect 79943 8336 80009 8359
rect 80095 8336 80177 8359
rect 80263 8336 80329 8359
rect 79943 8296 79952 8336
rect 79992 8296 80009 8336
rect 80095 8296 80116 8336
rect 80156 8296 80177 8336
rect 80263 8296 80280 8336
rect 80320 8296 80329 8336
rect 79943 8273 80009 8296
rect 80095 8273 80177 8296
rect 80263 8273 80329 8296
rect 79943 8254 80329 8273
rect 95063 8359 95449 8378
rect 95063 8336 95129 8359
rect 95215 8336 95297 8359
rect 95383 8336 95449 8359
rect 95063 8296 95072 8336
rect 95112 8296 95129 8336
rect 95215 8296 95236 8336
rect 95276 8296 95297 8336
rect 95383 8296 95400 8336
rect 95440 8296 95449 8336
rect 95063 8273 95129 8296
rect 95215 8273 95297 8296
rect 95383 8273 95449 8296
rect 95063 8254 95449 8273
rect 3103 7603 3489 7622
rect 3103 7580 3169 7603
rect 3255 7580 3337 7603
rect 3423 7580 3489 7603
rect 3103 7540 3112 7580
rect 3152 7540 3169 7580
rect 3255 7540 3276 7580
rect 3316 7540 3337 7580
rect 3423 7540 3440 7580
rect 3480 7540 3489 7580
rect 3103 7517 3169 7540
rect 3255 7517 3337 7540
rect 3423 7517 3489 7540
rect 3103 7498 3489 7517
rect 18223 7603 18609 7622
rect 18223 7580 18289 7603
rect 18375 7580 18457 7603
rect 18543 7580 18609 7603
rect 18223 7540 18232 7580
rect 18272 7540 18289 7580
rect 18375 7540 18396 7580
rect 18436 7540 18457 7580
rect 18543 7540 18560 7580
rect 18600 7540 18609 7580
rect 18223 7517 18289 7540
rect 18375 7517 18457 7540
rect 18543 7517 18609 7540
rect 18223 7498 18609 7517
rect 33343 7603 33729 7622
rect 33343 7580 33409 7603
rect 33495 7580 33577 7603
rect 33663 7580 33729 7603
rect 33343 7540 33352 7580
rect 33392 7540 33409 7580
rect 33495 7540 33516 7580
rect 33556 7540 33577 7580
rect 33663 7540 33680 7580
rect 33720 7540 33729 7580
rect 33343 7517 33409 7540
rect 33495 7517 33577 7540
rect 33663 7517 33729 7540
rect 33343 7498 33729 7517
rect 48463 7603 48849 7622
rect 48463 7580 48529 7603
rect 48615 7580 48697 7603
rect 48783 7580 48849 7603
rect 48463 7540 48472 7580
rect 48512 7540 48529 7580
rect 48615 7540 48636 7580
rect 48676 7540 48697 7580
rect 48783 7540 48800 7580
rect 48840 7540 48849 7580
rect 48463 7517 48529 7540
rect 48615 7517 48697 7540
rect 48783 7517 48849 7540
rect 48463 7498 48849 7517
rect 63583 7603 63969 7622
rect 63583 7580 63649 7603
rect 63735 7580 63817 7603
rect 63903 7580 63969 7603
rect 63583 7540 63592 7580
rect 63632 7540 63649 7580
rect 63735 7540 63756 7580
rect 63796 7540 63817 7580
rect 63903 7540 63920 7580
rect 63960 7540 63969 7580
rect 63583 7517 63649 7540
rect 63735 7517 63817 7540
rect 63903 7517 63969 7540
rect 63583 7498 63969 7517
rect 78703 7603 79089 7622
rect 78703 7580 78769 7603
rect 78855 7580 78937 7603
rect 79023 7580 79089 7603
rect 78703 7540 78712 7580
rect 78752 7540 78769 7580
rect 78855 7540 78876 7580
rect 78916 7540 78937 7580
rect 79023 7540 79040 7580
rect 79080 7540 79089 7580
rect 78703 7517 78769 7540
rect 78855 7517 78937 7540
rect 79023 7517 79089 7540
rect 78703 7498 79089 7517
rect 93823 7603 94209 7622
rect 93823 7580 93889 7603
rect 93975 7580 94057 7603
rect 94143 7580 94209 7603
rect 93823 7540 93832 7580
rect 93872 7540 93889 7580
rect 93975 7540 93996 7580
rect 94036 7540 94057 7580
rect 94143 7540 94160 7580
rect 94200 7540 94209 7580
rect 93823 7517 93889 7540
rect 93975 7517 94057 7540
rect 94143 7517 94209 7540
rect 93823 7498 94209 7517
rect 4343 6847 4729 6866
rect 4343 6824 4409 6847
rect 4495 6824 4577 6847
rect 4663 6824 4729 6847
rect 4343 6784 4352 6824
rect 4392 6784 4409 6824
rect 4495 6784 4516 6824
rect 4556 6784 4577 6824
rect 4663 6784 4680 6824
rect 4720 6784 4729 6824
rect 4343 6761 4409 6784
rect 4495 6761 4577 6784
rect 4663 6761 4729 6784
rect 4343 6742 4729 6761
rect 19463 6847 19849 6866
rect 19463 6824 19529 6847
rect 19615 6824 19697 6847
rect 19783 6824 19849 6847
rect 19463 6784 19472 6824
rect 19512 6784 19529 6824
rect 19615 6784 19636 6824
rect 19676 6784 19697 6824
rect 19783 6784 19800 6824
rect 19840 6784 19849 6824
rect 19463 6761 19529 6784
rect 19615 6761 19697 6784
rect 19783 6761 19849 6784
rect 19463 6742 19849 6761
rect 34583 6847 34969 6866
rect 34583 6824 34649 6847
rect 34735 6824 34817 6847
rect 34903 6824 34969 6847
rect 34583 6784 34592 6824
rect 34632 6784 34649 6824
rect 34735 6784 34756 6824
rect 34796 6784 34817 6824
rect 34903 6784 34920 6824
rect 34960 6784 34969 6824
rect 34583 6761 34649 6784
rect 34735 6761 34817 6784
rect 34903 6761 34969 6784
rect 34583 6742 34969 6761
rect 49703 6847 50089 6866
rect 49703 6824 49769 6847
rect 49855 6824 49937 6847
rect 50023 6824 50089 6847
rect 49703 6784 49712 6824
rect 49752 6784 49769 6824
rect 49855 6784 49876 6824
rect 49916 6784 49937 6824
rect 50023 6784 50040 6824
rect 50080 6784 50089 6824
rect 49703 6761 49769 6784
rect 49855 6761 49937 6784
rect 50023 6761 50089 6784
rect 49703 6742 50089 6761
rect 64823 6847 65209 6866
rect 64823 6824 64889 6847
rect 64975 6824 65057 6847
rect 65143 6824 65209 6847
rect 64823 6784 64832 6824
rect 64872 6784 64889 6824
rect 64975 6784 64996 6824
rect 65036 6784 65057 6824
rect 65143 6784 65160 6824
rect 65200 6784 65209 6824
rect 64823 6761 64889 6784
rect 64975 6761 65057 6784
rect 65143 6761 65209 6784
rect 64823 6742 65209 6761
rect 79943 6847 80329 6866
rect 79943 6824 80009 6847
rect 80095 6824 80177 6847
rect 80263 6824 80329 6847
rect 79943 6784 79952 6824
rect 79992 6784 80009 6824
rect 80095 6784 80116 6824
rect 80156 6784 80177 6824
rect 80263 6784 80280 6824
rect 80320 6784 80329 6824
rect 79943 6761 80009 6784
rect 80095 6761 80177 6784
rect 80263 6761 80329 6784
rect 79943 6742 80329 6761
rect 95063 6847 95449 6866
rect 95063 6824 95129 6847
rect 95215 6824 95297 6847
rect 95383 6824 95449 6847
rect 95063 6784 95072 6824
rect 95112 6784 95129 6824
rect 95215 6784 95236 6824
rect 95276 6784 95297 6824
rect 95383 6784 95400 6824
rect 95440 6784 95449 6824
rect 95063 6761 95129 6784
rect 95215 6761 95297 6784
rect 95383 6761 95449 6784
rect 95063 6742 95449 6761
rect 3103 6091 3489 6110
rect 3103 6068 3169 6091
rect 3255 6068 3337 6091
rect 3423 6068 3489 6091
rect 3103 6028 3112 6068
rect 3152 6028 3169 6068
rect 3255 6028 3276 6068
rect 3316 6028 3337 6068
rect 3423 6028 3440 6068
rect 3480 6028 3489 6068
rect 3103 6005 3169 6028
rect 3255 6005 3337 6028
rect 3423 6005 3489 6028
rect 3103 5986 3489 6005
rect 18223 6091 18609 6110
rect 18223 6068 18289 6091
rect 18375 6068 18457 6091
rect 18543 6068 18609 6091
rect 18223 6028 18232 6068
rect 18272 6028 18289 6068
rect 18375 6028 18396 6068
rect 18436 6028 18457 6068
rect 18543 6028 18560 6068
rect 18600 6028 18609 6068
rect 18223 6005 18289 6028
rect 18375 6005 18457 6028
rect 18543 6005 18609 6028
rect 18223 5986 18609 6005
rect 33343 6091 33729 6110
rect 33343 6068 33409 6091
rect 33495 6068 33577 6091
rect 33663 6068 33729 6091
rect 33343 6028 33352 6068
rect 33392 6028 33409 6068
rect 33495 6028 33516 6068
rect 33556 6028 33577 6068
rect 33663 6028 33680 6068
rect 33720 6028 33729 6068
rect 33343 6005 33409 6028
rect 33495 6005 33577 6028
rect 33663 6005 33729 6028
rect 33343 5986 33729 6005
rect 48463 6091 48849 6110
rect 48463 6068 48529 6091
rect 48615 6068 48697 6091
rect 48783 6068 48849 6091
rect 48463 6028 48472 6068
rect 48512 6028 48529 6068
rect 48615 6028 48636 6068
rect 48676 6028 48697 6068
rect 48783 6028 48800 6068
rect 48840 6028 48849 6068
rect 48463 6005 48529 6028
rect 48615 6005 48697 6028
rect 48783 6005 48849 6028
rect 48463 5986 48849 6005
rect 63583 6091 63969 6110
rect 63583 6068 63649 6091
rect 63735 6068 63817 6091
rect 63903 6068 63969 6091
rect 63583 6028 63592 6068
rect 63632 6028 63649 6068
rect 63735 6028 63756 6068
rect 63796 6028 63817 6068
rect 63903 6028 63920 6068
rect 63960 6028 63969 6068
rect 63583 6005 63649 6028
rect 63735 6005 63817 6028
rect 63903 6005 63969 6028
rect 63583 5986 63969 6005
rect 78703 6091 79089 6110
rect 78703 6068 78769 6091
rect 78855 6068 78937 6091
rect 79023 6068 79089 6091
rect 78703 6028 78712 6068
rect 78752 6028 78769 6068
rect 78855 6028 78876 6068
rect 78916 6028 78937 6068
rect 79023 6028 79040 6068
rect 79080 6028 79089 6068
rect 78703 6005 78769 6028
rect 78855 6005 78937 6028
rect 79023 6005 79089 6028
rect 78703 5986 79089 6005
rect 93823 6091 94209 6110
rect 93823 6068 93889 6091
rect 93975 6068 94057 6091
rect 94143 6068 94209 6091
rect 93823 6028 93832 6068
rect 93872 6028 93889 6068
rect 93975 6028 93996 6068
rect 94036 6028 94057 6068
rect 94143 6028 94160 6068
rect 94200 6028 94209 6068
rect 93823 6005 93889 6028
rect 93975 6005 94057 6028
rect 94143 6005 94209 6028
rect 93823 5986 94209 6005
rect 4343 5335 4729 5354
rect 4343 5312 4409 5335
rect 4495 5312 4577 5335
rect 4663 5312 4729 5335
rect 4343 5272 4352 5312
rect 4392 5272 4409 5312
rect 4495 5272 4516 5312
rect 4556 5272 4577 5312
rect 4663 5272 4680 5312
rect 4720 5272 4729 5312
rect 4343 5249 4409 5272
rect 4495 5249 4577 5272
rect 4663 5249 4729 5272
rect 4343 5230 4729 5249
rect 19463 5335 19849 5354
rect 19463 5312 19529 5335
rect 19615 5312 19697 5335
rect 19783 5312 19849 5335
rect 19463 5272 19472 5312
rect 19512 5272 19529 5312
rect 19615 5272 19636 5312
rect 19676 5272 19697 5312
rect 19783 5272 19800 5312
rect 19840 5272 19849 5312
rect 19463 5249 19529 5272
rect 19615 5249 19697 5272
rect 19783 5249 19849 5272
rect 19463 5230 19849 5249
rect 34583 5335 34969 5354
rect 34583 5312 34649 5335
rect 34735 5312 34817 5335
rect 34903 5312 34969 5335
rect 34583 5272 34592 5312
rect 34632 5272 34649 5312
rect 34735 5272 34756 5312
rect 34796 5272 34817 5312
rect 34903 5272 34920 5312
rect 34960 5272 34969 5312
rect 34583 5249 34649 5272
rect 34735 5249 34817 5272
rect 34903 5249 34969 5272
rect 34583 5230 34969 5249
rect 49703 5335 50089 5354
rect 49703 5312 49769 5335
rect 49855 5312 49937 5335
rect 50023 5312 50089 5335
rect 49703 5272 49712 5312
rect 49752 5272 49769 5312
rect 49855 5272 49876 5312
rect 49916 5272 49937 5312
rect 50023 5272 50040 5312
rect 50080 5272 50089 5312
rect 49703 5249 49769 5272
rect 49855 5249 49937 5272
rect 50023 5249 50089 5272
rect 49703 5230 50089 5249
rect 64823 5335 65209 5354
rect 64823 5312 64889 5335
rect 64975 5312 65057 5335
rect 65143 5312 65209 5335
rect 64823 5272 64832 5312
rect 64872 5272 64889 5312
rect 64975 5272 64996 5312
rect 65036 5272 65057 5312
rect 65143 5272 65160 5312
rect 65200 5272 65209 5312
rect 64823 5249 64889 5272
rect 64975 5249 65057 5272
rect 65143 5249 65209 5272
rect 64823 5230 65209 5249
rect 79943 5335 80329 5354
rect 79943 5312 80009 5335
rect 80095 5312 80177 5335
rect 80263 5312 80329 5335
rect 79943 5272 79952 5312
rect 79992 5272 80009 5312
rect 80095 5272 80116 5312
rect 80156 5272 80177 5312
rect 80263 5272 80280 5312
rect 80320 5272 80329 5312
rect 79943 5249 80009 5272
rect 80095 5249 80177 5272
rect 80263 5249 80329 5272
rect 79943 5230 80329 5249
rect 95063 5335 95449 5354
rect 95063 5312 95129 5335
rect 95215 5312 95297 5335
rect 95383 5312 95449 5335
rect 95063 5272 95072 5312
rect 95112 5272 95129 5312
rect 95215 5272 95236 5312
rect 95276 5272 95297 5312
rect 95383 5272 95400 5312
rect 95440 5272 95449 5312
rect 95063 5249 95129 5272
rect 95215 5249 95297 5272
rect 95383 5249 95449 5272
rect 95063 5230 95449 5249
rect 3103 4579 3489 4598
rect 3103 4556 3169 4579
rect 3255 4556 3337 4579
rect 3423 4556 3489 4579
rect 3103 4516 3112 4556
rect 3152 4516 3169 4556
rect 3255 4516 3276 4556
rect 3316 4516 3337 4556
rect 3423 4516 3440 4556
rect 3480 4516 3489 4556
rect 3103 4493 3169 4516
rect 3255 4493 3337 4516
rect 3423 4493 3489 4516
rect 3103 4474 3489 4493
rect 18223 4579 18609 4598
rect 18223 4556 18289 4579
rect 18375 4556 18457 4579
rect 18543 4556 18609 4579
rect 18223 4516 18232 4556
rect 18272 4516 18289 4556
rect 18375 4516 18396 4556
rect 18436 4516 18457 4556
rect 18543 4516 18560 4556
rect 18600 4516 18609 4556
rect 18223 4493 18289 4516
rect 18375 4493 18457 4516
rect 18543 4493 18609 4516
rect 18223 4474 18609 4493
rect 33343 4579 33729 4598
rect 33343 4556 33409 4579
rect 33495 4556 33577 4579
rect 33663 4556 33729 4579
rect 33343 4516 33352 4556
rect 33392 4516 33409 4556
rect 33495 4516 33516 4556
rect 33556 4516 33577 4556
rect 33663 4516 33680 4556
rect 33720 4516 33729 4556
rect 33343 4493 33409 4516
rect 33495 4493 33577 4516
rect 33663 4493 33729 4516
rect 33343 4474 33729 4493
rect 48463 4579 48849 4598
rect 48463 4556 48529 4579
rect 48615 4556 48697 4579
rect 48783 4556 48849 4579
rect 48463 4516 48472 4556
rect 48512 4516 48529 4556
rect 48615 4516 48636 4556
rect 48676 4516 48697 4556
rect 48783 4516 48800 4556
rect 48840 4516 48849 4556
rect 48463 4493 48529 4516
rect 48615 4493 48697 4516
rect 48783 4493 48849 4516
rect 48463 4474 48849 4493
rect 63583 4579 63969 4598
rect 63583 4556 63649 4579
rect 63735 4556 63817 4579
rect 63903 4556 63969 4579
rect 63583 4516 63592 4556
rect 63632 4516 63649 4556
rect 63735 4516 63756 4556
rect 63796 4516 63817 4556
rect 63903 4516 63920 4556
rect 63960 4516 63969 4556
rect 63583 4493 63649 4516
rect 63735 4493 63817 4516
rect 63903 4493 63969 4516
rect 63583 4474 63969 4493
rect 78703 4579 79089 4598
rect 78703 4556 78769 4579
rect 78855 4556 78937 4579
rect 79023 4556 79089 4579
rect 78703 4516 78712 4556
rect 78752 4516 78769 4556
rect 78855 4516 78876 4556
rect 78916 4516 78937 4556
rect 79023 4516 79040 4556
rect 79080 4516 79089 4556
rect 78703 4493 78769 4516
rect 78855 4493 78937 4516
rect 79023 4493 79089 4516
rect 78703 4474 79089 4493
rect 93823 4579 94209 4598
rect 93823 4556 93889 4579
rect 93975 4556 94057 4579
rect 94143 4556 94209 4579
rect 93823 4516 93832 4556
rect 93872 4516 93889 4556
rect 93975 4516 93996 4556
rect 94036 4516 94057 4556
rect 94143 4516 94160 4556
rect 94200 4516 94209 4556
rect 93823 4493 93889 4516
rect 93975 4493 94057 4516
rect 94143 4493 94209 4516
rect 93823 4474 94209 4493
rect 4343 3823 4729 3842
rect 4343 3800 4409 3823
rect 4495 3800 4577 3823
rect 4663 3800 4729 3823
rect 4343 3760 4352 3800
rect 4392 3760 4409 3800
rect 4495 3760 4516 3800
rect 4556 3760 4577 3800
rect 4663 3760 4680 3800
rect 4720 3760 4729 3800
rect 4343 3737 4409 3760
rect 4495 3737 4577 3760
rect 4663 3737 4729 3760
rect 4343 3718 4729 3737
rect 19463 3823 19849 3842
rect 19463 3800 19529 3823
rect 19615 3800 19697 3823
rect 19783 3800 19849 3823
rect 19463 3760 19472 3800
rect 19512 3760 19529 3800
rect 19615 3760 19636 3800
rect 19676 3760 19697 3800
rect 19783 3760 19800 3800
rect 19840 3760 19849 3800
rect 19463 3737 19529 3760
rect 19615 3737 19697 3760
rect 19783 3737 19849 3760
rect 19463 3718 19849 3737
rect 34583 3823 34969 3842
rect 34583 3800 34649 3823
rect 34735 3800 34817 3823
rect 34903 3800 34969 3823
rect 34583 3760 34592 3800
rect 34632 3760 34649 3800
rect 34735 3760 34756 3800
rect 34796 3760 34817 3800
rect 34903 3760 34920 3800
rect 34960 3760 34969 3800
rect 34583 3737 34649 3760
rect 34735 3737 34817 3760
rect 34903 3737 34969 3760
rect 34583 3718 34969 3737
rect 49703 3823 50089 3842
rect 49703 3800 49769 3823
rect 49855 3800 49937 3823
rect 50023 3800 50089 3823
rect 49703 3760 49712 3800
rect 49752 3760 49769 3800
rect 49855 3760 49876 3800
rect 49916 3760 49937 3800
rect 50023 3760 50040 3800
rect 50080 3760 50089 3800
rect 49703 3737 49769 3760
rect 49855 3737 49937 3760
rect 50023 3737 50089 3760
rect 49703 3718 50089 3737
rect 64823 3823 65209 3842
rect 64823 3800 64889 3823
rect 64975 3800 65057 3823
rect 65143 3800 65209 3823
rect 64823 3760 64832 3800
rect 64872 3760 64889 3800
rect 64975 3760 64996 3800
rect 65036 3760 65057 3800
rect 65143 3760 65160 3800
rect 65200 3760 65209 3800
rect 64823 3737 64889 3760
rect 64975 3737 65057 3760
rect 65143 3737 65209 3760
rect 64823 3718 65209 3737
rect 79943 3823 80329 3842
rect 79943 3800 80009 3823
rect 80095 3800 80177 3823
rect 80263 3800 80329 3823
rect 79943 3760 79952 3800
rect 79992 3760 80009 3800
rect 80095 3760 80116 3800
rect 80156 3760 80177 3800
rect 80263 3760 80280 3800
rect 80320 3760 80329 3800
rect 79943 3737 80009 3760
rect 80095 3737 80177 3760
rect 80263 3737 80329 3760
rect 79943 3718 80329 3737
rect 95063 3823 95449 3842
rect 95063 3800 95129 3823
rect 95215 3800 95297 3823
rect 95383 3800 95449 3823
rect 95063 3760 95072 3800
rect 95112 3760 95129 3800
rect 95215 3760 95236 3800
rect 95276 3760 95297 3800
rect 95383 3760 95400 3800
rect 95440 3760 95449 3800
rect 95063 3737 95129 3760
rect 95215 3737 95297 3760
rect 95383 3737 95449 3760
rect 95063 3718 95449 3737
rect 3103 3067 3489 3086
rect 3103 3044 3169 3067
rect 3255 3044 3337 3067
rect 3423 3044 3489 3067
rect 3103 3004 3112 3044
rect 3152 3004 3169 3044
rect 3255 3004 3276 3044
rect 3316 3004 3337 3044
rect 3423 3004 3440 3044
rect 3480 3004 3489 3044
rect 3103 2981 3169 3004
rect 3255 2981 3337 3004
rect 3423 2981 3489 3004
rect 3103 2962 3489 2981
rect 18223 3067 18609 3086
rect 18223 3044 18289 3067
rect 18375 3044 18457 3067
rect 18543 3044 18609 3067
rect 18223 3004 18232 3044
rect 18272 3004 18289 3044
rect 18375 3004 18396 3044
rect 18436 3004 18457 3044
rect 18543 3004 18560 3044
rect 18600 3004 18609 3044
rect 18223 2981 18289 3004
rect 18375 2981 18457 3004
rect 18543 2981 18609 3004
rect 18223 2962 18609 2981
rect 33343 3067 33729 3086
rect 33343 3044 33409 3067
rect 33495 3044 33577 3067
rect 33663 3044 33729 3067
rect 33343 3004 33352 3044
rect 33392 3004 33409 3044
rect 33495 3004 33516 3044
rect 33556 3004 33577 3044
rect 33663 3004 33680 3044
rect 33720 3004 33729 3044
rect 33343 2981 33409 3004
rect 33495 2981 33577 3004
rect 33663 2981 33729 3004
rect 33343 2962 33729 2981
rect 48463 3067 48849 3086
rect 48463 3044 48529 3067
rect 48615 3044 48697 3067
rect 48783 3044 48849 3067
rect 48463 3004 48472 3044
rect 48512 3004 48529 3044
rect 48615 3004 48636 3044
rect 48676 3004 48697 3044
rect 48783 3004 48800 3044
rect 48840 3004 48849 3044
rect 48463 2981 48529 3004
rect 48615 2981 48697 3004
rect 48783 2981 48849 3004
rect 48463 2962 48849 2981
rect 63583 3067 63969 3086
rect 63583 3044 63649 3067
rect 63735 3044 63817 3067
rect 63903 3044 63969 3067
rect 63583 3004 63592 3044
rect 63632 3004 63649 3044
rect 63735 3004 63756 3044
rect 63796 3004 63817 3044
rect 63903 3004 63920 3044
rect 63960 3004 63969 3044
rect 63583 2981 63649 3004
rect 63735 2981 63817 3004
rect 63903 2981 63969 3004
rect 63583 2962 63969 2981
rect 78703 3067 79089 3086
rect 78703 3044 78769 3067
rect 78855 3044 78937 3067
rect 79023 3044 79089 3067
rect 78703 3004 78712 3044
rect 78752 3004 78769 3044
rect 78855 3004 78876 3044
rect 78916 3004 78937 3044
rect 79023 3004 79040 3044
rect 79080 3004 79089 3044
rect 78703 2981 78769 3004
rect 78855 2981 78937 3004
rect 79023 2981 79089 3004
rect 78703 2962 79089 2981
rect 93823 3067 94209 3086
rect 93823 3044 93889 3067
rect 93975 3044 94057 3067
rect 94143 3044 94209 3067
rect 93823 3004 93832 3044
rect 93872 3004 93889 3044
rect 93975 3004 93996 3044
rect 94036 3004 94057 3044
rect 94143 3004 94160 3044
rect 94200 3004 94209 3044
rect 93823 2981 93889 3004
rect 93975 2981 94057 3004
rect 94143 2981 94209 3004
rect 93823 2962 94209 2981
rect 4343 2311 4729 2330
rect 4343 2288 4409 2311
rect 4495 2288 4577 2311
rect 4663 2288 4729 2311
rect 4343 2248 4352 2288
rect 4392 2248 4409 2288
rect 4495 2248 4516 2288
rect 4556 2248 4577 2288
rect 4663 2248 4680 2288
rect 4720 2248 4729 2288
rect 4343 2225 4409 2248
rect 4495 2225 4577 2248
rect 4663 2225 4729 2248
rect 4343 2206 4729 2225
rect 19463 2311 19849 2330
rect 19463 2288 19529 2311
rect 19615 2288 19697 2311
rect 19783 2288 19849 2311
rect 19463 2248 19472 2288
rect 19512 2248 19529 2288
rect 19615 2248 19636 2288
rect 19676 2248 19697 2288
rect 19783 2248 19800 2288
rect 19840 2248 19849 2288
rect 19463 2225 19529 2248
rect 19615 2225 19697 2248
rect 19783 2225 19849 2248
rect 19463 2206 19849 2225
rect 34583 2311 34969 2330
rect 34583 2288 34649 2311
rect 34735 2288 34817 2311
rect 34903 2288 34969 2311
rect 34583 2248 34592 2288
rect 34632 2248 34649 2288
rect 34735 2248 34756 2288
rect 34796 2248 34817 2288
rect 34903 2248 34920 2288
rect 34960 2248 34969 2288
rect 34583 2225 34649 2248
rect 34735 2225 34817 2248
rect 34903 2225 34969 2248
rect 34583 2206 34969 2225
rect 49703 2311 50089 2330
rect 49703 2288 49769 2311
rect 49855 2288 49937 2311
rect 50023 2288 50089 2311
rect 49703 2248 49712 2288
rect 49752 2248 49769 2288
rect 49855 2248 49876 2288
rect 49916 2248 49937 2288
rect 50023 2248 50040 2288
rect 50080 2248 50089 2288
rect 49703 2225 49769 2248
rect 49855 2225 49937 2248
rect 50023 2225 50089 2248
rect 49703 2206 50089 2225
rect 64823 2311 65209 2330
rect 64823 2288 64889 2311
rect 64975 2288 65057 2311
rect 65143 2288 65209 2311
rect 64823 2248 64832 2288
rect 64872 2248 64889 2288
rect 64975 2248 64996 2288
rect 65036 2248 65057 2288
rect 65143 2248 65160 2288
rect 65200 2248 65209 2288
rect 64823 2225 64889 2248
rect 64975 2225 65057 2248
rect 65143 2225 65209 2248
rect 64823 2206 65209 2225
rect 79943 2311 80329 2330
rect 79943 2288 80009 2311
rect 80095 2288 80177 2311
rect 80263 2288 80329 2311
rect 79943 2248 79952 2288
rect 79992 2248 80009 2288
rect 80095 2248 80116 2288
rect 80156 2248 80177 2288
rect 80263 2248 80280 2288
rect 80320 2248 80329 2288
rect 79943 2225 80009 2248
rect 80095 2225 80177 2248
rect 80263 2225 80329 2248
rect 79943 2206 80329 2225
rect 95063 2311 95449 2330
rect 95063 2288 95129 2311
rect 95215 2288 95297 2311
rect 95383 2288 95449 2311
rect 95063 2248 95072 2288
rect 95112 2248 95129 2288
rect 95215 2248 95236 2288
rect 95276 2248 95297 2288
rect 95383 2248 95400 2288
rect 95440 2248 95449 2288
rect 95063 2225 95129 2248
rect 95215 2225 95297 2248
rect 95383 2225 95449 2248
rect 95063 2206 95449 2225
rect 3103 1555 3489 1574
rect 3103 1532 3169 1555
rect 3255 1532 3337 1555
rect 3423 1532 3489 1555
rect 3103 1492 3112 1532
rect 3152 1492 3169 1532
rect 3255 1492 3276 1532
rect 3316 1492 3337 1532
rect 3423 1492 3440 1532
rect 3480 1492 3489 1532
rect 3103 1469 3169 1492
rect 3255 1469 3337 1492
rect 3423 1469 3489 1492
rect 3103 1450 3489 1469
rect 18223 1555 18609 1574
rect 18223 1532 18289 1555
rect 18375 1532 18457 1555
rect 18543 1532 18609 1555
rect 18223 1492 18232 1532
rect 18272 1492 18289 1532
rect 18375 1492 18396 1532
rect 18436 1492 18457 1532
rect 18543 1492 18560 1532
rect 18600 1492 18609 1532
rect 18223 1469 18289 1492
rect 18375 1469 18457 1492
rect 18543 1469 18609 1492
rect 18223 1450 18609 1469
rect 33343 1555 33729 1574
rect 33343 1532 33409 1555
rect 33495 1532 33577 1555
rect 33663 1532 33729 1555
rect 33343 1492 33352 1532
rect 33392 1492 33409 1532
rect 33495 1492 33516 1532
rect 33556 1492 33577 1532
rect 33663 1492 33680 1532
rect 33720 1492 33729 1532
rect 33343 1469 33409 1492
rect 33495 1469 33577 1492
rect 33663 1469 33729 1492
rect 33343 1450 33729 1469
rect 48463 1555 48849 1574
rect 48463 1532 48529 1555
rect 48615 1532 48697 1555
rect 48783 1532 48849 1555
rect 48463 1492 48472 1532
rect 48512 1492 48529 1532
rect 48615 1492 48636 1532
rect 48676 1492 48697 1532
rect 48783 1492 48800 1532
rect 48840 1492 48849 1532
rect 48463 1469 48529 1492
rect 48615 1469 48697 1492
rect 48783 1469 48849 1492
rect 48463 1450 48849 1469
rect 63583 1555 63969 1574
rect 63583 1532 63649 1555
rect 63735 1532 63817 1555
rect 63903 1532 63969 1555
rect 63583 1492 63592 1532
rect 63632 1492 63649 1532
rect 63735 1492 63756 1532
rect 63796 1492 63817 1532
rect 63903 1492 63920 1532
rect 63960 1492 63969 1532
rect 63583 1469 63649 1492
rect 63735 1469 63817 1492
rect 63903 1469 63969 1492
rect 63583 1450 63969 1469
rect 78703 1555 79089 1574
rect 78703 1532 78769 1555
rect 78855 1532 78937 1555
rect 79023 1532 79089 1555
rect 78703 1492 78712 1532
rect 78752 1492 78769 1532
rect 78855 1492 78876 1532
rect 78916 1492 78937 1532
rect 79023 1492 79040 1532
rect 79080 1492 79089 1532
rect 78703 1469 78769 1492
rect 78855 1469 78937 1492
rect 79023 1469 79089 1492
rect 78703 1450 79089 1469
rect 93823 1555 94209 1574
rect 93823 1532 93889 1555
rect 93975 1532 94057 1555
rect 94143 1532 94209 1555
rect 93823 1492 93832 1532
rect 93872 1492 93889 1532
rect 93975 1492 93996 1532
rect 94036 1492 94057 1532
rect 94143 1492 94160 1532
rect 94200 1492 94209 1532
rect 93823 1469 93889 1492
rect 93975 1469 94057 1492
rect 94143 1469 94209 1492
rect 93823 1450 94209 1469
rect 4343 799 4729 818
rect 4343 776 4409 799
rect 4495 776 4577 799
rect 4663 776 4729 799
rect 4343 736 4352 776
rect 4392 736 4409 776
rect 4495 736 4516 776
rect 4556 736 4577 776
rect 4663 736 4680 776
rect 4720 736 4729 776
rect 4343 713 4409 736
rect 4495 713 4577 736
rect 4663 713 4729 736
rect 4343 694 4729 713
rect 19463 799 19849 818
rect 19463 776 19529 799
rect 19615 776 19697 799
rect 19783 776 19849 799
rect 19463 736 19472 776
rect 19512 736 19529 776
rect 19615 736 19636 776
rect 19676 736 19697 776
rect 19783 736 19800 776
rect 19840 736 19849 776
rect 19463 713 19529 736
rect 19615 713 19697 736
rect 19783 713 19849 736
rect 19463 694 19849 713
rect 34583 799 34969 818
rect 34583 776 34649 799
rect 34735 776 34817 799
rect 34903 776 34969 799
rect 34583 736 34592 776
rect 34632 736 34649 776
rect 34735 736 34756 776
rect 34796 736 34817 776
rect 34903 736 34920 776
rect 34960 736 34969 776
rect 34583 713 34649 736
rect 34735 713 34817 736
rect 34903 713 34969 736
rect 34583 694 34969 713
rect 49703 799 50089 818
rect 49703 776 49769 799
rect 49855 776 49937 799
rect 50023 776 50089 799
rect 49703 736 49712 776
rect 49752 736 49769 776
rect 49855 736 49876 776
rect 49916 736 49937 776
rect 50023 736 50040 776
rect 50080 736 50089 776
rect 49703 713 49769 736
rect 49855 713 49937 736
rect 50023 713 50089 736
rect 49703 694 50089 713
rect 64823 799 65209 818
rect 64823 776 64889 799
rect 64975 776 65057 799
rect 65143 776 65209 799
rect 64823 736 64832 776
rect 64872 736 64889 776
rect 64975 736 64996 776
rect 65036 736 65057 776
rect 65143 736 65160 776
rect 65200 736 65209 776
rect 64823 713 64889 736
rect 64975 713 65057 736
rect 65143 713 65209 736
rect 64823 694 65209 713
rect 79943 799 80329 818
rect 79943 776 80009 799
rect 80095 776 80177 799
rect 80263 776 80329 799
rect 79943 736 79952 776
rect 79992 736 80009 776
rect 80095 736 80116 776
rect 80156 736 80177 776
rect 80263 736 80280 776
rect 80320 736 80329 776
rect 79943 713 80009 736
rect 80095 713 80177 736
rect 80263 713 80329 736
rect 79943 694 80329 713
rect 95063 799 95449 818
rect 95063 776 95129 799
rect 95215 776 95297 799
rect 95383 776 95449 799
rect 95063 736 95072 776
rect 95112 736 95129 776
rect 95215 736 95236 776
rect 95276 736 95297 776
rect 95383 736 95400 776
rect 95440 736 95449 776
rect 95063 713 95129 736
rect 95215 713 95297 736
rect 95383 713 95449 736
rect 95063 694 95449 713
<< via5 >>
rect 4409 38576 4495 38599
rect 4577 38576 4663 38599
rect 4409 38536 4434 38576
rect 4434 38536 4474 38576
rect 4474 38536 4495 38576
rect 4577 38536 4598 38576
rect 4598 38536 4638 38576
rect 4638 38536 4663 38576
rect 4409 38513 4495 38536
rect 4577 38513 4663 38536
rect 19529 38576 19615 38599
rect 19697 38576 19783 38599
rect 19529 38536 19554 38576
rect 19554 38536 19594 38576
rect 19594 38536 19615 38576
rect 19697 38536 19718 38576
rect 19718 38536 19758 38576
rect 19758 38536 19783 38576
rect 19529 38513 19615 38536
rect 19697 38513 19783 38536
rect 34649 38576 34735 38599
rect 34817 38576 34903 38599
rect 34649 38536 34674 38576
rect 34674 38536 34714 38576
rect 34714 38536 34735 38576
rect 34817 38536 34838 38576
rect 34838 38536 34878 38576
rect 34878 38536 34903 38576
rect 34649 38513 34735 38536
rect 34817 38513 34903 38536
rect 49769 38576 49855 38599
rect 49937 38576 50023 38599
rect 49769 38536 49794 38576
rect 49794 38536 49834 38576
rect 49834 38536 49855 38576
rect 49937 38536 49958 38576
rect 49958 38536 49998 38576
rect 49998 38536 50023 38576
rect 49769 38513 49855 38536
rect 49937 38513 50023 38536
rect 64889 38576 64975 38599
rect 65057 38576 65143 38599
rect 64889 38536 64914 38576
rect 64914 38536 64954 38576
rect 64954 38536 64975 38576
rect 65057 38536 65078 38576
rect 65078 38536 65118 38576
rect 65118 38536 65143 38576
rect 64889 38513 64975 38536
rect 65057 38513 65143 38536
rect 80009 38576 80095 38599
rect 80177 38576 80263 38599
rect 80009 38536 80034 38576
rect 80034 38536 80074 38576
rect 80074 38536 80095 38576
rect 80177 38536 80198 38576
rect 80198 38536 80238 38576
rect 80238 38536 80263 38576
rect 80009 38513 80095 38536
rect 80177 38513 80263 38536
rect 95129 38576 95215 38599
rect 95297 38576 95383 38599
rect 95129 38536 95154 38576
rect 95154 38536 95194 38576
rect 95194 38536 95215 38576
rect 95297 38536 95318 38576
rect 95318 38536 95358 38576
rect 95358 38536 95383 38576
rect 95129 38513 95215 38536
rect 95297 38513 95383 38536
rect 3169 37820 3255 37843
rect 3337 37820 3423 37843
rect 3169 37780 3194 37820
rect 3194 37780 3234 37820
rect 3234 37780 3255 37820
rect 3337 37780 3358 37820
rect 3358 37780 3398 37820
rect 3398 37780 3423 37820
rect 3169 37757 3255 37780
rect 3337 37757 3423 37780
rect 18289 37820 18375 37843
rect 18457 37820 18543 37843
rect 18289 37780 18314 37820
rect 18314 37780 18354 37820
rect 18354 37780 18375 37820
rect 18457 37780 18478 37820
rect 18478 37780 18518 37820
rect 18518 37780 18543 37820
rect 18289 37757 18375 37780
rect 18457 37757 18543 37780
rect 33409 37820 33495 37843
rect 33577 37820 33663 37843
rect 33409 37780 33434 37820
rect 33434 37780 33474 37820
rect 33474 37780 33495 37820
rect 33577 37780 33598 37820
rect 33598 37780 33638 37820
rect 33638 37780 33663 37820
rect 33409 37757 33495 37780
rect 33577 37757 33663 37780
rect 48529 37820 48615 37843
rect 48697 37820 48783 37843
rect 48529 37780 48554 37820
rect 48554 37780 48594 37820
rect 48594 37780 48615 37820
rect 48697 37780 48718 37820
rect 48718 37780 48758 37820
rect 48758 37780 48783 37820
rect 48529 37757 48615 37780
rect 48697 37757 48783 37780
rect 63649 37820 63735 37843
rect 63817 37820 63903 37843
rect 63649 37780 63674 37820
rect 63674 37780 63714 37820
rect 63714 37780 63735 37820
rect 63817 37780 63838 37820
rect 63838 37780 63878 37820
rect 63878 37780 63903 37820
rect 63649 37757 63735 37780
rect 63817 37757 63903 37780
rect 78769 37820 78855 37843
rect 78937 37820 79023 37843
rect 78769 37780 78794 37820
rect 78794 37780 78834 37820
rect 78834 37780 78855 37820
rect 78937 37780 78958 37820
rect 78958 37780 78998 37820
rect 78998 37780 79023 37820
rect 78769 37757 78855 37780
rect 78937 37757 79023 37780
rect 93889 37820 93975 37843
rect 94057 37820 94143 37843
rect 93889 37780 93914 37820
rect 93914 37780 93954 37820
rect 93954 37780 93975 37820
rect 94057 37780 94078 37820
rect 94078 37780 94118 37820
rect 94118 37780 94143 37820
rect 93889 37757 93975 37780
rect 94057 37757 94143 37780
rect 4409 37064 4495 37087
rect 4577 37064 4663 37087
rect 4409 37024 4434 37064
rect 4434 37024 4474 37064
rect 4474 37024 4495 37064
rect 4577 37024 4598 37064
rect 4598 37024 4638 37064
rect 4638 37024 4663 37064
rect 4409 37001 4495 37024
rect 4577 37001 4663 37024
rect 19529 37064 19615 37087
rect 19697 37064 19783 37087
rect 19529 37024 19554 37064
rect 19554 37024 19594 37064
rect 19594 37024 19615 37064
rect 19697 37024 19718 37064
rect 19718 37024 19758 37064
rect 19758 37024 19783 37064
rect 19529 37001 19615 37024
rect 19697 37001 19783 37024
rect 34649 37064 34735 37087
rect 34817 37064 34903 37087
rect 34649 37024 34674 37064
rect 34674 37024 34714 37064
rect 34714 37024 34735 37064
rect 34817 37024 34838 37064
rect 34838 37024 34878 37064
rect 34878 37024 34903 37064
rect 34649 37001 34735 37024
rect 34817 37001 34903 37024
rect 49769 37064 49855 37087
rect 49937 37064 50023 37087
rect 49769 37024 49794 37064
rect 49794 37024 49834 37064
rect 49834 37024 49855 37064
rect 49937 37024 49958 37064
rect 49958 37024 49998 37064
rect 49998 37024 50023 37064
rect 49769 37001 49855 37024
rect 49937 37001 50023 37024
rect 64889 37064 64975 37087
rect 65057 37064 65143 37087
rect 64889 37024 64914 37064
rect 64914 37024 64954 37064
rect 64954 37024 64975 37064
rect 65057 37024 65078 37064
rect 65078 37024 65118 37064
rect 65118 37024 65143 37064
rect 64889 37001 64975 37024
rect 65057 37001 65143 37024
rect 80009 37064 80095 37087
rect 80177 37064 80263 37087
rect 80009 37024 80034 37064
rect 80034 37024 80074 37064
rect 80074 37024 80095 37064
rect 80177 37024 80198 37064
rect 80198 37024 80238 37064
rect 80238 37024 80263 37064
rect 80009 37001 80095 37024
rect 80177 37001 80263 37024
rect 95129 37064 95215 37087
rect 95297 37064 95383 37087
rect 95129 37024 95154 37064
rect 95154 37024 95194 37064
rect 95194 37024 95215 37064
rect 95297 37024 95318 37064
rect 95318 37024 95358 37064
rect 95358 37024 95383 37064
rect 95129 37001 95215 37024
rect 95297 37001 95383 37024
rect 3169 36308 3255 36331
rect 3337 36308 3423 36331
rect 3169 36268 3194 36308
rect 3194 36268 3234 36308
rect 3234 36268 3255 36308
rect 3337 36268 3358 36308
rect 3358 36268 3398 36308
rect 3398 36268 3423 36308
rect 3169 36245 3255 36268
rect 3337 36245 3423 36268
rect 18289 36308 18375 36331
rect 18457 36308 18543 36331
rect 18289 36268 18314 36308
rect 18314 36268 18354 36308
rect 18354 36268 18375 36308
rect 18457 36268 18478 36308
rect 18478 36268 18518 36308
rect 18518 36268 18543 36308
rect 18289 36245 18375 36268
rect 18457 36245 18543 36268
rect 33409 36308 33495 36331
rect 33577 36308 33663 36331
rect 33409 36268 33434 36308
rect 33434 36268 33474 36308
rect 33474 36268 33495 36308
rect 33577 36268 33598 36308
rect 33598 36268 33638 36308
rect 33638 36268 33663 36308
rect 33409 36245 33495 36268
rect 33577 36245 33663 36268
rect 48529 36308 48615 36331
rect 48697 36308 48783 36331
rect 48529 36268 48554 36308
rect 48554 36268 48594 36308
rect 48594 36268 48615 36308
rect 48697 36268 48718 36308
rect 48718 36268 48758 36308
rect 48758 36268 48783 36308
rect 48529 36245 48615 36268
rect 48697 36245 48783 36268
rect 63649 36308 63735 36331
rect 63817 36308 63903 36331
rect 63649 36268 63674 36308
rect 63674 36268 63714 36308
rect 63714 36268 63735 36308
rect 63817 36268 63838 36308
rect 63838 36268 63878 36308
rect 63878 36268 63903 36308
rect 63649 36245 63735 36268
rect 63817 36245 63903 36268
rect 78769 36308 78855 36331
rect 78937 36308 79023 36331
rect 78769 36268 78794 36308
rect 78794 36268 78834 36308
rect 78834 36268 78855 36308
rect 78937 36268 78958 36308
rect 78958 36268 78998 36308
rect 78998 36268 79023 36308
rect 78769 36245 78855 36268
rect 78937 36245 79023 36268
rect 93889 36308 93975 36331
rect 94057 36308 94143 36331
rect 93889 36268 93914 36308
rect 93914 36268 93954 36308
rect 93954 36268 93975 36308
rect 94057 36268 94078 36308
rect 94078 36268 94118 36308
rect 94118 36268 94143 36308
rect 93889 36245 93975 36268
rect 94057 36245 94143 36268
rect 4409 35552 4495 35575
rect 4577 35552 4663 35575
rect 4409 35512 4434 35552
rect 4434 35512 4474 35552
rect 4474 35512 4495 35552
rect 4577 35512 4598 35552
rect 4598 35512 4638 35552
rect 4638 35512 4663 35552
rect 4409 35489 4495 35512
rect 4577 35489 4663 35512
rect 19529 35552 19615 35575
rect 19697 35552 19783 35575
rect 19529 35512 19554 35552
rect 19554 35512 19594 35552
rect 19594 35512 19615 35552
rect 19697 35512 19718 35552
rect 19718 35512 19758 35552
rect 19758 35512 19783 35552
rect 19529 35489 19615 35512
rect 19697 35489 19783 35512
rect 34649 35552 34735 35575
rect 34817 35552 34903 35575
rect 34649 35512 34674 35552
rect 34674 35512 34714 35552
rect 34714 35512 34735 35552
rect 34817 35512 34838 35552
rect 34838 35512 34878 35552
rect 34878 35512 34903 35552
rect 34649 35489 34735 35512
rect 34817 35489 34903 35512
rect 49769 35552 49855 35575
rect 49937 35552 50023 35575
rect 49769 35512 49794 35552
rect 49794 35512 49834 35552
rect 49834 35512 49855 35552
rect 49937 35512 49958 35552
rect 49958 35512 49998 35552
rect 49998 35512 50023 35552
rect 49769 35489 49855 35512
rect 49937 35489 50023 35512
rect 64889 35552 64975 35575
rect 65057 35552 65143 35575
rect 64889 35512 64914 35552
rect 64914 35512 64954 35552
rect 64954 35512 64975 35552
rect 65057 35512 65078 35552
rect 65078 35512 65118 35552
rect 65118 35512 65143 35552
rect 64889 35489 64975 35512
rect 65057 35489 65143 35512
rect 80009 35552 80095 35575
rect 80177 35552 80263 35575
rect 80009 35512 80034 35552
rect 80034 35512 80074 35552
rect 80074 35512 80095 35552
rect 80177 35512 80198 35552
rect 80198 35512 80238 35552
rect 80238 35512 80263 35552
rect 80009 35489 80095 35512
rect 80177 35489 80263 35512
rect 95129 35552 95215 35575
rect 95297 35552 95383 35575
rect 95129 35512 95154 35552
rect 95154 35512 95194 35552
rect 95194 35512 95215 35552
rect 95297 35512 95318 35552
rect 95318 35512 95358 35552
rect 95358 35512 95383 35552
rect 95129 35489 95215 35512
rect 95297 35489 95383 35512
rect 3169 34796 3255 34819
rect 3337 34796 3423 34819
rect 3169 34756 3194 34796
rect 3194 34756 3234 34796
rect 3234 34756 3255 34796
rect 3337 34756 3358 34796
rect 3358 34756 3398 34796
rect 3398 34756 3423 34796
rect 3169 34733 3255 34756
rect 3337 34733 3423 34756
rect 18289 34796 18375 34819
rect 18457 34796 18543 34819
rect 18289 34756 18314 34796
rect 18314 34756 18354 34796
rect 18354 34756 18375 34796
rect 18457 34756 18478 34796
rect 18478 34756 18518 34796
rect 18518 34756 18543 34796
rect 18289 34733 18375 34756
rect 18457 34733 18543 34756
rect 33409 34796 33495 34819
rect 33577 34796 33663 34819
rect 33409 34756 33434 34796
rect 33434 34756 33474 34796
rect 33474 34756 33495 34796
rect 33577 34756 33598 34796
rect 33598 34756 33638 34796
rect 33638 34756 33663 34796
rect 33409 34733 33495 34756
rect 33577 34733 33663 34756
rect 48529 34796 48615 34819
rect 48697 34796 48783 34819
rect 48529 34756 48554 34796
rect 48554 34756 48594 34796
rect 48594 34756 48615 34796
rect 48697 34756 48718 34796
rect 48718 34756 48758 34796
rect 48758 34756 48783 34796
rect 48529 34733 48615 34756
rect 48697 34733 48783 34756
rect 63649 34796 63735 34819
rect 63817 34796 63903 34819
rect 63649 34756 63674 34796
rect 63674 34756 63714 34796
rect 63714 34756 63735 34796
rect 63817 34756 63838 34796
rect 63838 34756 63878 34796
rect 63878 34756 63903 34796
rect 63649 34733 63735 34756
rect 63817 34733 63903 34756
rect 78769 34796 78855 34819
rect 78937 34796 79023 34819
rect 78769 34756 78794 34796
rect 78794 34756 78834 34796
rect 78834 34756 78855 34796
rect 78937 34756 78958 34796
rect 78958 34756 78998 34796
rect 78998 34756 79023 34796
rect 78769 34733 78855 34756
rect 78937 34733 79023 34756
rect 93889 34796 93975 34819
rect 94057 34796 94143 34819
rect 93889 34756 93914 34796
rect 93914 34756 93954 34796
rect 93954 34756 93975 34796
rect 94057 34756 94078 34796
rect 94078 34756 94118 34796
rect 94118 34756 94143 34796
rect 93889 34733 93975 34756
rect 94057 34733 94143 34756
rect 4409 34040 4495 34063
rect 4577 34040 4663 34063
rect 4409 34000 4434 34040
rect 4434 34000 4474 34040
rect 4474 34000 4495 34040
rect 4577 34000 4598 34040
rect 4598 34000 4638 34040
rect 4638 34000 4663 34040
rect 4409 33977 4495 34000
rect 4577 33977 4663 34000
rect 19529 34040 19615 34063
rect 19697 34040 19783 34063
rect 19529 34000 19554 34040
rect 19554 34000 19594 34040
rect 19594 34000 19615 34040
rect 19697 34000 19718 34040
rect 19718 34000 19758 34040
rect 19758 34000 19783 34040
rect 19529 33977 19615 34000
rect 19697 33977 19783 34000
rect 34649 34040 34735 34063
rect 34817 34040 34903 34063
rect 34649 34000 34674 34040
rect 34674 34000 34714 34040
rect 34714 34000 34735 34040
rect 34817 34000 34838 34040
rect 34838 34000 34878 34040
rect 34878 34000 34903 34040
rect 34649 33977 34735 34000
rect 34817 33977 34903 34000
rect 49769 34040 49855 34063
rect 49937 34040 50023 34063
rect 49769 34000 49794 34040
rect 49794 34000 49834 34040
rect 49834 34000 49855 34040
rect 49937 34000 49958 34040
rect 49958 34000 49998 34040
rect 49998 34000 50023 34040
rect 49769 33977 49855 34000
rect 49937 33977 50023 34000
rect 64889 34040 64975 34063
rect 65057 34040 65143 34063
rect 64889 34000 64914 34040
rect 64914 34000 64954 34040
rect 64954 34000 64975 34040
rect 65057 34000 65078 34040
rect 65078 34000 65118 34040
rect 65118 34000 65143 34040
rect 64889 33977 64975 34000
rect 65057 33977 65143 34000
rect 80009 34040 80095 34063
rect 80177 34040 80263 34063
rect 80009 34000 80034 34040
rect 80034 34000 80074 34040
rect 80074 34000 80095 34040
rect 80177 34000 80198 34040
rect 80198 34000 80238 34040
rect 80238 34000 80263 34040
rect 80009 33977 80095 34000
rect 80177 33977 80263 34000
rect 95129 34040 95215 34063
rect 95297 34040 95383 34063
rect 95129 34000 95154 34040
rect 95154 34000 95194 34040
rect 95194 34000 95215 34040
rect 95297 34000 95318 34040
rect 95318 34000 95358 34040
rect 95358 34000 95383 34040
rect 95129 33977 95215 34000
rect 95297 33977 95383 34000
rect 3169 33284 3255 33307
rect 3337 33284 3423 33307
rect 3169 33244 3194 33284
rect 3194 33244 3234 33284
rect 3234 33244 3255 33284
rect 3337 33244 3358 33284
rect 3358 33244 3398 33284
rect 3398 33244 3423 33284
rect 3169 33221 3255 33244
rect 3337 33221 3423 33244
rect 18289 33284 18375 33307
rect 18457 33284 18543 33307
rect 18289 33244 18314 33284
rect 18314 33244 18354 33284
rect 18354 33244 18375 33284
rect 18457 33244 18478 33284
rect 18478 33244 18518 33284
rect 18518 33244 18543 33284
rect 18289 33221 18375 33244
rect 18457 33221 18543 33244
rect 33409 33284 33495 33307
rect 33577 33284 33663 33307
rect 33409 33244 33434 33284
rect 33434 33244 33474 33284
rect 33474 33244 33495 33284
rect 33577 33244 33598 33284
rect 33598 33244 33638 33284
rect 33638 33244 33663 33284
rect 33409 33221 33495 33244
rect 33577 33221 33663 33244
rect 48529 33284 48615 33307
rect 48697 33284 48783 33307
rect 48529 33244 48554 33284
rect 48554 33244 48594 33284
rect 48594 33244 48615 33284
rect 48697 33244 48718 33284
rect 48718 33244 48758 33284
rect 48758 33244 48783 33284
rect 48529 33221 48615 33244
rect 48697 33221 48783 33244
rect 63649 33284 63735 33307
rect 63817 33284 63903 33307
rect 63649 33244 63674 33284
rect 63674 33244 63714 33284
rect 63714 33244 63735 33284
rect 63817 33244 63838 33284
rect 63838 33244 63878 33284
rect 63878 33244 63903 33284
rect 63649 33221 63735 33244
rect 63817 33221 63903 33244
rect 78769 33284 78855 33307
rect 78937 33284 79023 33307
rect 78769 33244 78794 33284
rect 78794 33244 78834 33284
rect 78834 33244 78855 33284
rect 78937 33244 78958 33284
rect 78958 33244 78998 33284
rect 78998 33244 79023 33284
rect 78769 33221 78855 33244
rect 78937 33221 79023 33244
rect 93889 33284 93975 33307
rect 94057 33284 94143 33307
rect 93889 33244 93914 33284
rect 93914 33244 93954 33284
rect 93954 33244 93975 33284
rect 94057 33244 94078 33284
rect 94078 33244 94118 33284
rect 94118 33244 94143 33284
rect 93889 33221 93975 33244
rect 94057 33221 94143 33244
rect 4409 32528 4495 32551
rect 4577 32528 4663 32551
rect 4409 32488 4434 32528
rect 4434 32488 4474 32528
rect 4474 32488 4495 32528
rect 4577 32488 4598 32528
rect 4598 32488 4638 32528
rect 4638 32488 4663 32528
rect 4409 32465 4495 32488
rect 4577 32465 4663 32488
rect 19529 32528 19615 32551
rect 19697 32528 19783 32551
rect 19529 32488 19554 32528
rect 19554 32488 19594 32528
rect 19594 32488 19615 32528
rect 19697 32488 19718 32528
rect 19718 32488 19758 32528
rect 19758 32488 19783 32528
rect 19529 32465 19615 32488
rect 19697 32465 19783 32488
rect 34649 32528 34735 32551
rect 34817 32528 34903 32551
rect 34649 32488 34674 32528
rect 34674 32488 34714 32528
rect 34714 32488 34735 32528
rect 34817 32488 34838 32528
rect 34838 32488 34878 32528
rect 34878 32488 34903 32528
rect 34649 32465 34735 32488
rect 34817 32465 34903 32488
rect 49769 32528 49855 32551
rect 49937 32528 50023 32551
rect 49769 32488 49794 32528
rect 49794 32488 49834 32528
rect 49834 32488 49855 32528
rect 49937 32488 49958 32528
rect 49958 32488 49998 32528
rect 49998 32488 50023 32528
rect 49769 32465 49855 32488
rect 49937 32465 50023 32488
rect 64889 32528 64975 32551
rect 65057 32528 65143 32551
rect 64889 32488 64914 32528
rect 64914 32488 64954 32528
rect 64954 32488 64975 32528
rect 65057 32488 65078 32528
rect 65078 32488 65118 32528
rect 65118 32488 65143 32528
rect 64889 32465 64975 32488
rect 65057 32465 65143 32488
rect 80009 32528 80095 32551
rect 80177 32528 80263 32551
rect 80009 32488 80034 32528
rect 80034 32488 80074 32528
rect 80074 32488 80095 32528
rect 80177 32488 80198 32528
rect 80198 32488 80238 32528
rect 80238 32488 80263 32528
rect 80009 32465 80095 32488
rect 80177 32465 80263 32488
rect 95129 32528 95215 32551
rect 95297 32528 95383 32551
rect 95129 32488 95154 32528
rect 95154 32488 95194 32528
rect 95194 32488 95215 32528
rect 95297 32488 95318 32528
rect 95318 32488 95358 32528
rect 95358 32488 95383 32528
rect 95129 32465 95215 32488
rect 95297 32465 95383 32488
rect 3169 31772 3255 31795
rect 3337 31772 3423 31795
rect 3169 31732 3194 31772
rect 3194 31732 3234 31772
rect 3234 31732 3255 31772
rect 3337 31732 3358 31772
rect 3358 31732 3398 31772
rect 3398 31732 3423 31772
rect 3169 31709 3255 31732
rect 3337 31709 3423 31732
rect 18289 31772 18375 31795
rect 18457 31772 18543 31795
rect 18289 31732 18314 31772
rect 18314 31732 18354 31772
rect 18354 31732 18375 31772
rect 18457 31732 18478 31772
rect 18478 31732 18518 31772
rect 18518 31732 18543 31772
rect 18289 31709 18375 31732
rect 18457 31709 18543 31732
rect 33409 31772 33495 31795
rect 33577 31772 33663 31795
rect 33409 31732 33434 31772
rect 33434 31732 33474 31772
rect 33474 31732 33495 31772
rect 33577 31732 33598 31772
rect 33598 31732 33638 31772
rect 33638 31732 33663 31772
rect 33409 31709 33495 31732
rect 33577 31709 33663 31732
rect 48529 31772 48615 31795
rect 48697 31772 48783 31795
rect 48529 31732 48554 31772
rect 48554 31732 48594 31772
rect 48594 31732 48615 31772
rect 48697 31732 48718 31772
rect 48718 31732 48758 31772
rect 48758 31732 48783 31772
rect 48529 31709 48615 31732
rect 48697 31709 48783 31732
rect 63649 31772 63735 31795
rect 63817 31772 63903 31795
rect 63649 31732 63674 31772
rect 63674 31732 63714 31772
rect 63714 31732 63735 31772
rect 63817 31732 63838 31772
rect 63838 31732 63878 31772
rect 63878 31732 63903 31772
rect 63649 31709 63735 31732
rect 63817 31709 63903 31732
rect 78769 31772 78855 31795
rect 78937 31772 79023 31795
rect 78769 31732 78794 31772
rect 78794 31732 78834 31772
rect 78834 31732 78855 31772
rect 78937 31732 78958 31772
rect 78958 31732 78998 31772
rect 78998 31732 79023 31772
rect 78769 31709 78855 31732
rect 78937 31709 79023 31732
rect 93889 31772 93975 31795
rect 94057 31772 94143 31795
rect 93889 31732 93914 31772
rect 93914 31732 93954 31772
rect 93954 31732 93975 31772
rect 94057 31732 94078 31772
rect 94078 31732 94118 31772
rect 94118 31732 94143 31772
rect 93889 31709 93975 31732
rect 94057 31709 94143 31732
rect 4409 31016 4495 31039
rect 4577 31016 4663 31039
rect 4409 30976 4434 31016
rect 4434 30976 4474 31016
rect 4474 30976 4495 31016
rect 4577 30976 4598 31016
rect 4598 30976 4638 31016
rect 4638 30976 4663 31016
rect 4409 30953 4495 30976
rect 4577 30953 4663 30976
rect 19529 31016 19615 31039
rect 19697 31016 19783 31039
rect 19529 30976 19554 31016
rect 19554 30976 19594 31016
rect 19594 30976 19615 31016
rect 19697 30976 19718 31016
rect 19718 30976 19758 31016
rect 19758 30976 19783 31016
rect 19529 30953 19615 30976
rect 19697 30953 19783 30976
rect 34649 31016 34735 31039
rect 34817 31016 34903 31039
rect 34649 30976 34674 31016
rect 34674 30976 34714 31016
rect 34714 30976 34735 31016
rect 34817 30976 34838 31016
rect 34838 30976 34878 31016
rect 34878 30976 34903 31016
rect 34649 30953 34735 30976
rect 34817 30953 34903 30976
rect 49769 31016 49855 31039
rect 49937 31016 50023 31039
rect 49769 30976 49794 31016
rect 49794 30976 49834 31016
rect 49834 30976 49855 31016
rect 49937 30976 49958 31016
rect 49958 30976 49998 31016
rect 49998 30976 50023 31016
rect 49769 30953 49855 30976
rect 49937 30953 50023 30976
rect 64889 31016 64975 31039
rect 65057 31016 65143 31039
rect 64889 30976 64914 31016
rect 64914 30976 64954 31016
rect 64954 30976 64975 31016
rect 65057 30976 65078 31016
rect 65078 30976 65118 31016
rect 65118 30976 65143 31016
rect 64889 30953 64975 30976
rect 65057 30953 65143 30976
rect 80009 31016 80095 31039
rect 80177 31016 80263 31039
rect 80009 30976 80034 31016
rect 80034 30976 80074 31016
rect 80074 30976 80095 31016
rect 80177 30976 80198 31016
rect 80198 30976 80238 31016
rect 80238 30976 80263 31016
rect 80009 30953 80095 30976
rect 80177 30953 80263 30976
rect 95129 31016 95215 31039
rect 95297 31016 95383 31039
rect 95129 30976 95154 31016
rect 95154 30976 95194 31016
rect 95194 30976 95215 31016
rect 95297 30976 95318 31016
rect 95318 30976 95358 31016
rect 95358 30976 95383 31016
rect 95129 30953 95215 30976
rect 95297 30953 95383 30976
rect 3169 30260 3255 30283
rect 3337 30260 3423 30283
rect 3169 30220 3194 30260
rect 3194 30220 3234 30260
rect 3234 30220 3255 30260
rect 3337 30220 3358 30260
rect 3358 30220 3398 30260
rect 3398 30220 3423 30260
rect 3169 30197 3255 30220
rect 3337 30197 3423 30220
rect 18289 30260 18375 30283
rect 18457 30260 18543 30283
rect 18289 30220 18314 30260
rect 18314 30220 18354 30260
rect 18354 30220 18375 30260
rect 18457 30220 18478 30260
rect 18478 30220 18518 30260
rect 18518 30220 18543 30260
rect 18289 30197 18375 30220
rect 18457 30197 18543 30220
rect 33409 30260 33495 30283
rect 33577 30260 33663 30283
rect 33409 30220 33434 30260
rect 33434 30220 33474 30260
rect 33474 30220 33495 30260
rect 33577 30220 33598 30260
rect 33598 30220 33638 30260
rect 33638 30220 33663 30260
rect 33409 30197 33495 30220
rect 33577 30197 33663 30220
rect 48529 30260 48615 30283
rect 48697 30260 48783 30283
rect 48529 30220 48554 30260
rect 48554 30220 48594 30260
rect 48594 30220 48615 30260
rect 48697 30220 48718 30260
rect 48718 30220 48758 30260
rect 48758 30220 48783 30260
rect 48529 30197 48615 30220
rect 48697 30197 48783 30220
rect 63649 30260 63735 30283
rect 63817 30260 63903 30283
rect 63649 30220 63674 30260
rect 63674 30220 63714 30260
rect 63714 30220 63735 30260
rect 63817 30220 63838 30260
rect 63838 30220 63878 30260
rect 63878 30220 63903 30260
rect 63649 30197 63735 30220
rect 63817 30197 63903 30220
rect 78769 30260 78855 30283
rect 78937 30260 79023 30283
rect 78769 30220 78794 30260
rect 78794 30220 78834 30260
rect 78834 30220 78855 30260
rect 78937 30220 78958 30260
rect 78958 30220 78998 30260
rect 78998 30220 79023 30260
rect 78769 30197 78855 30220
rect 78937 30197 79023 30220
rect 93889 30260 93975 30283
rect 94057 30260 94143 30283
rect 93889 30220 93914 30260
rect 93914 30220 93954 30260
rect 93954 30220 93975 30260
rect 94057 30220 94078 30260
rect 94078 30220 94118 30260
rect 94118 30220 94143 30260
rect 93889 30197 93975 30220
rect 94057 30197 94143 30220
rect 4409 29504 4495 29527
rect 4577 29504 4663 29527
rect 4409 29464 4434 29504
rect 4434 29464 4474 29504
rect 4474 29464 4495 29504
rect 4577 29464 4598 29504
rect 4598 29464 4638 29504
rect 4638 29464 4663 29504
rect 4409 29441 4495 29464
rect 4577 29441 4663 29464
rect 19529 29504 19615 29527
rect 19697 29504 19783 29527
rect 19529 29464 19554 29504
rect 19554 29464 19594 29504
rect 19594 29464 19615 29504
rect 19697 29464 19718 29504
rect 19718 29464 19758 29504
rect 19758 29464 19783 29504
rect 19529 29441 19615 29464
rect 19697 29441 19783 29464
rect 34649 29504 34735 29527
rect 34817 29504 34903 29527
rect 34649 29464 34674 29504
rect 34674 29464 34714 29504
rect 34714 29464 34735 29504
rect 34817 29464 34838 29504
rect 34838 29464 34878 29504
rect 34878 29464 34903 29504
rect 34649 29441 34735 29464
rect 34817 29441 34903 29464
rect 49769 29504 49855 29527
rect 49937 29504 50023 29527
rect 49769 29464 49794 29504
rect 49794 29464 49834 29504
rect 49834 29464 49855 29504
rect 49937 29464 49958 29504
rect 49958 29464 49998 29504
rect 49998 29464 50023 29504
rect 49769 29441 49855 29464
rect 49937 29441 50023 29464
rect 64889 29504 64975 29527
rect 65057 29504 65143 29527
rect 64889 29464 64914 29504
rect 64914 29464 64954 29504
rect 64954 29464 64975 29504
rect 65057 29464 65078 29504
rect 65078 29464 65118 29504
rect 65118 29464 65143 29504
rect 64889 29441 64975 29464
rect 65057 29441 65143 29464
rect 80009 29504 80095 29527
rect 80177 29504 80263 29527
rect 80009 29464 80034 29504
rect 80034 29464 80074 29504
rect 80074 29464 80095 29504
rect 80177 29464 80198 29504
rect 80198 29464 80238 29504
rect 80238 29464 80263 29504
rect 80009 29441 80095 29464
rect 80177 29441 80263 29464
rect 95129 29504 95215 29527
rect 95297 29504 95383 29527
rect 95129 29464 95154 29504
rect 95154 29464 95194 29504
rect 95194 29464 95215 29504
rect 95297 29464 95318 29504
rect 95318 29464 95358 29504
rect 95358 29464 95383 29504
rect 95129 29441 95215 29464
rect 95297 29441 95383 29464
rect 3169 28748 3255 28771
rect 3337 28748 3423 28771
rect 3169 28708 3194 28748
rect 3194 28708 3234 28748
rect 3234 28708 3255 28748
rect 3337 28708 3358 28748
rect 3358 28708 3398 28748
rect 3398 28708 3423 28748
rect 3169 28685 3255 28708
rect 3337 28685 3423 28708
rect 18289 28748 18375 28771
rect 18457 28748 18543 28771
rect 18289 28708 18314 28748
rect 18314 28708 18354 28748
rect 18354 28708 18375 28748
rect 18457 28708 18478 28748
rect 18478 28708 18518 28748
rect 18518 28708 18543 28748
rect 18289 28685 18375 28708
rect 18457 28685 18543 28708
rect 33409 28748 33495 28771
rect 33577 28748 33663 28771
rect 33409 28708 33434 28748
rect 33434 28708 33474 28748
rect 33474 28708 33495 28748
rect 33577 28708 33598 28748
rect 33598 28708 33638 28748
rect 33638 28708 33663 28748
rect 33409 28685 33495 28708
rect 33577 28685 33663 28708
rect 48529 28748 48615 28771
rect 48697 28748 48783 28771
rect 48529 28708 48554 28748
rect 48554 28708 48594 28748
rect 48594 28708 48615 28748
rect 48697 28708 48718 28748
rect 48718 28708 48758 28748
rect 48758 28708 48783 28748
rect 48529 28685 48615 28708
rect 48697 28685 48783 28708
rect 63649 28748 63735 28771
rect 63817 28748 63903 28771
rect 63649 28708 63674 28748
rect 63674 28708 63714 28748
rect 63714 28708 63735 28748
rect 63817 28708 63838 28748
rect 63838 28708 63878 28748
rect 63878 28708 63903 28748
rect 63649 28685 63735 28708
rect 63817 28685 63903 28708
rect 78769 28748 78855 28771
rect 78937 28748 79023 28771
rect 78769 28708 78794 28748
rect 78794 28708 78834 28748
rect 78834 28708 78855 28748
rect 78937 28708 78958 28748
rect 78958 28708 78998 28748
rect 78998 28708 79023 28748
rect 78769 28685 78855 28708
rect 78937 28685 79023 28708
rect 93889 28748 93975 28771
rect 94057 28748 94143 28771
rect 93889 28708 93914 28748
rect 93914 28708 93954 28748
rect 93954 28708 93975 28748
rect 94057 28708 94078 28748
rect 94078 28708 94118 28748
rect 94118 28708 94143 28748
rect 93889 28685 93975 28708
rect 94057 28685 94143 28708
rect 4409 27992 4495 28015
rect 4577 27992 4663 28015
rect 4409 27952 4434 27992
rect 4434 27952 4474 27992
rect 4474 27952 4495 27992
rect 4577 27952 4598 27992
rect 4598 27952 4638 27992
rect 4638 27952 4663 27992
rect 4409 27929 4495 27952
rect 4577 27929 4663 27952
rect 19529 27992 19615 28015
rect 19697 27992 19783 28015
rect 19529 27952 19554 27992
rect 19554 27952 19594 27992
rect 19594 27952 19615 27992
rect 19697 27952 19718 27992
rect 19718 27952 19758 27992
rect 19758 27952 19783 27992
rect 19529 27929 19615 27952
rect 19697 27929 19783 27952
rect 34649 27992 34735 28015
rect 34817 27992 34903 28015
rect 34649 27952 34674 27992
rect 34674 27952 34714 27992
rect 34714 27952 34735 27992
rect 34817 27952 34838 27992
rect 34838 27952 34878 27992
rect 34878 27952 34903 27992
rect 34649 27929 34735 27952
rect 34817 27929 34903 27952
rect 49769 27992 49855 28015
rect 49937 27992 50023 28015
rect 49769 27952 49794 27992
rect 49794 27952 49834 27992
rect 49834 27952 49855 27992
rect 49937 27952 49958 27992
rect 49958 27952 49998 27992
rect 49998 27952 50023 27992
rect 49769 27929 49855 27952
rect 49937 27929 50023 27952
rect 64889 27992 64975 28015
rect 65057 27992 65143 28015
rect 64889 27952 64914 27992
rect 64914 27952 64954 27992
rect 64954 27952 64975 27992
rect 65057 27952 65078 27992
rect 65078 27952 65118 27992
rect 65118 27952 65143 27992
rect 64889 27929 64975 27952
rect 65057 27929 65143 27952
rect 80009 27992 80095 28015
rect 80177 27992 80263 28015
rect 80009 27952 80034 27992
rect 80034 27952 80074 27992
rect 80074 27952 80095 27992
rect 80177 27952 80198 27992
rect 80198 27952 80238 27992
rect 80238 27952 80263 27992
rect 80009 27929 80095 27952
rect 80177 27929 80263 27952
rect 95129 27992 95215 28015
rect 95297 27992 95383 28015
rect 95129 27952 95154 27992
rect 95154 27952 95194 27992
rect 95194 27952 95215 27992
rect 95297 27952 95318 27992
rect 95318 27952 95358 27992
rect 95358 27952 95383 27992
rect 95129 27929 95215 27952
rect 95297 27929 95383 27952
rect 3169 27236 3255 27259
rect 3337 27236 3423 27259
rect 3169 27196 3194 27236
rect 3194 27196 3234 27236
rect 3234 27196 3255 27236
rect 3337 27196 3358 27236
rect 3358 27196 3398 27236
rect 3398 27196 3423 27236
rect 3169 27173 3255 27196
rect 3337 27173 3423 27196
rect 18289 27236 18375 27259
rect 18457 27236 18543 27259
rect 18289 27196 18314 27236
rect 18314 27196 18354 27236
rect 18354 27196 18375 27236
rect 18457 27196 18478 27236
rect 18478 27196 18518 27236
rect 18518 27196 18543 27236
rect 18289 27173 18375 27196
rect 18457 27173 18543 27196
rect 33409 27236 33495 27259
rect 33577 27236 33663 27259
rect 33409 27196 33434 27236
rect 33434 27196 33474 27236
rect 33474 27196 33495 27236
rect 33577 27196 33598 27236
rect 33598 27196 33638 27236
rect 33638 27196 33663 27236
rect 33409 27173 33495 27196
rect 33577 27173 33663 27196
rect 48529 27236 48615 27259
rect 48697 27236 48783 27259
rect 48529 27196 48554 27236
rect 48554 27196 48594 27236
rect 48594 27196 48615 27236
rect 48697 27196 48718 27236
rect 48718 27196 48758 27236
rect 48758 27196 48783 27236
rect 48529 27173 48615 27196
rect 48697 27173 48783 27196
rect 63649 27236 63735 27259
rect 63817 27236 63903 27259
rect 63649 27196 63674 27236
rect 63674 27196 63714 27236
rect 63714 27196 63735 27236
rect 63817 27196 63838 27236
rect 63838 27196 63878 27236
rect 63878 27196 63903 27236
rect 63649 27173 63735 27196
rect 63817 27173 63903 27196
rect 78769 27236 78855 27259
rect 78937 27236 79023 27259
rect 78769 27196 78794 27236
rect 78794 27196 78834 27236
rect 78834 27196 78855 27236
rect 78937 27196 78958 27236
rect 78958 27196 78998 27236
rect 78998 27196 79023 27236
rect 78769 27173 78855 27196
rect 78937 27173 79023 27196
rect 93889 27236 93975 27259
rect 94057 27236 94143 27259
rect 93889 27196 93914 27236
rect 93914 27196 93954 27236
rect 93954 27196 93975 27236
rect 94057 27196 94078 27236
rect 94078 27196 94118 27236
rect 94118 27196 94143 27236
rect 93889 27173 93975 27196
rect 94057 27173 94143 27196
rect 4409 26480 4495 26503
rect 4577 26480 4663 26503
rect 4409 26440 4434 26480
rect 4434 26440 4474 26480
rect 4474 26440 4495 26480
rect 4577 26440 4598 26480
rect 4598 26440 4638 26480
rect 4638 26440 4663 26480
rect 4409 26417 4495 26440
rect 4577 26417 4663 26440
rect 19529 26480 19615 26503
rect 19697 26480 19783 26503
rect 19529 26440 19554 26480
rect 19554 26440 19594 26480
rect 19594 26440 19615 26480
rect 19697 26440 19718 26480
rect 19718 26440 19758 26480
rect 19758 26440 19783 26480
rect 19529 26417 19615 26440
rect 19697 26417 19783 26440
rect 34649 26480 34735 26503
rect 34817 26480 34903 26503
rect 34649 26440 34674 26480
rect 34674 26440 34714 26480
rect 34714 26440 34735 26480
rect 34817 26440 34838 26480
rect 34838 26440 34878 26480
rect 34878 26440 34903 26480
rect 34649 26417 34735 26440
rect 34817 26417 34903 26440
rect 49769 26480 49855 26503
rect 49937 26480 50023 26503
rect 49769 26440 49794 26480
rect 49794 26440 49834 26480
rect 49834 26440 49855 26480
rect 49937 26440 49958 26480
rect 49958 26440 49998 26480
rect 49998 26440 50023 26480
rect 49769 26417 49855 26440
rect 49937 26417 50023 26440
rect 64889 26480 64975 26503
rect 65057 26480 65143 26503
rect 64889 26440 64914 26480
rect 64914 26440 64954 26480
rect 64954 26440 64975 26480
rect 65057 26440 65078 26480
rect 65078 26440 65118 26480
rect 65118 26440 65143 26480
rect 64889 26417 64975 26440
rect 65057 26417 65143 26440
rect 80009 26480 80095 26503
rect 80177 26480 80263 26503
rect 80009 26440 80034 26480
rect 80034 26440 80074 26480
rect 80074 26440 80095 26480
rect 80177 26440 80198 26480
rect 80198 26440 80238 26480
rect 80238 26440 80263 26480
rect 80009 26417 80095 26440
rect 80177 26417 80263 26440
rect 95129 26480 95215 26503
rect 95297 26480 95383 26503
rect 95129 26440 95154 26480
rect 95154 26440 95194 26480
rect 95194 26440 95215 26480
rect 95297 26440 95318 26480
rect 95318 26440 95358 26480
rect 95358 26440 95383 26480
rect 95129 26417 95215 26440
rect 95297 26417 95383 26440
rect 3169 25724 3255 25747
rect 3337 25724 3423 25747
rect 3169 25684 3194 25724
rect 3194 25684 3234 25724
rect 3234 25684 3255 25724
rect 3337 25684 3358 25724
rect 3358 25684 3398 25724
rect 3398 25684 3423 25724
rect 3169 25661 3255 25684
rect 3337 25661 3423 25684
rect 18289 25724 18375 25747
rect 18457 25724 18543 25747
rect 18289 25684 18314 25724
rect 18314 25684 18354 25724
rect 18354 25684 18375 25724
rect 18457 25684 18478 25724
rect 18478 25684 18518 25724
rect 18518 25684 18543 25724
rect 18289 25661 18375 25684
rect 18457 25661 18543 25684
rect 33409 25724 33495 25747
rect 33577 25724 33663 25747
rect 33409 25684 33434 25724
rect 33434 25684 33474 25724
rect 33474 25684 33495 25724
rect 33577 25684 33598 25724
rect 33598 25684 33638 25724
rect 33638 25684 33663 25724
rect 33409 25661 33495 25684
rect 33577 25661 33663 25684
rect 48529 25724 48615 25747
rect 48697 25724 48783 25747
rect 48529 25684 48554 25724
rect 48554 25684 48594 25724
rect 48594 25684 48615 25724
rect 48697 25684 48718 25724
rect 48718 25684 48758 25724
rect 48758 25684 48783 25724
rect 48529 25661 48615 25684
rect 48697 25661 48783 25684
rect 63649 25724 63735 25747
rect 63817 25724 63903 25747
rect 63649 25684 63674 25724
rect 63674 25684 63714 25724
rect 63714 25684 63735 25724
rect 63817 25684 63838 25724
rect 63838 25684 63878 25724
rect 63878 25684 63903 25724
rect 63649 25661 63735 25684
rect 63817 25661 63903 25684
rect 78769 25724 78855 25747
rect 78937 25724 79023 25747
rect 78769 25684 78794 25724
rect 78794 25684 78834 25724
rect 78834 25684 78855 25724
rect 78937 25684 78958 25724
rect 78958 25684 78998 25724
rect 78998 25684 79023 25724
rect 78769 25661 78855 25684
rect 78937 25661 79023 25684
rect 93889 25724 93975 25747
rect 94057 25724 94143 25747
rect 93889 25684 93914 25724
rect 93914 25684 93954 25724
rect 93954 25684 93975 25724
rect 94057 25684 94078 25724
rect 94078 25684 94118 25724
rect 94118 25684 94143 25724
rect 93889 25661 93975 25684
rect 94057 25661 94143 25684
rect 4409 24968 4495 24991
rect 4577 24968 4663 24991
rect 4409 24928 4434 24968
rect 4434 24928 4474 24968
rect 4474 24928 4495 24968
rect 4577 24928 4598 24968
rect 4598 24928 4638 24968
rect 4638 24928 4663 24968
rect 4409 24905 4495 24928
rect 4577 24905 4663 24928
rect 19529 24968 19615 24991
rect 19697 24968 19783 24991
rect 19529 24928 19554 24968
rect 19554 24928 19594 24968
rect 19594 24928 19615 24968
rect 19697 24928 19718 24968
rect 19718 24928 19758 24968
rect 19758 24928 19783 24968
rect 19529 24905 19615 24928
rect 19697 24905 19783 24928
rect 34649 24968 34735 24991
rect 34817 24968 34903 24991
rect 34649 24928 34674 24968
rect 34674 24928 34714 24968
rect 34714 24928 34735 24968
rect 34817 24928 34838 24968
rect 34838 24928 34878 24968
rect 34878 24928 34903 24968
rect 34649 24905 34735 24928
rect 34817 24905 34903 24928
rect 49769 24968 49855 24991
rect 49937 24968 50023 24991
rect 49769 24928 49794 24968
rect 49794 24928 49834 24968
rect 49834 24928 49855 24968
rect 49937 24928 49958 24968
rect 49958 24928 49998 24968
rect 49998 24928 50023 24968
rect 49769 24905 49855 24928
rect 49937 24905 50023 24928
rect 64889 24968 64975 24991
rect 65057 24968 65143 24991
rect 64889 24928 64914 24968
rect 64914 24928 64954 24968
rect 64954 24928 64975 24968
rect 65057 24928 65078 24968
rect 65078 24928 65118 24968
rect 65118 24928 65143 24968
rect 64889 24905 64975 24928
rect 65057 24905 65143 24928
rect 80009 24968 80095 24991
rect 80177 24968 80263 24991
rect 80009 24928 80034 24968
rect 80034 24928 80074 24968
rect 80074 24928 80095 24968
rect 80177 24928 80198 24968
rect 80198 24928 80238 24968
rect 80238 24928 80263 24968
rect 80009 24905 80095 24928
rect 80177 24905 80263 24928
rect 95129 24968 95215 24991
rect 95297 24968 95383 24991
rect 95129 24928 95154 24968
rect 95154 24928 95194 24968
rect 95194 24928 95215 24968
rect 95297 24928 95318 24968
rect 95318 24928 95358 24968
rect 95358 24928 95383 24968
rect 95129 24905 95215 24928
rect 95297 24905 95383 24928
rect 3169 24212 3255 24235
rect 3337 24212 3423 24235
rect 3169 24172 3194 24212
rect 3194 24172 3234 24212
rect 3234 24172 3255 24212
rect 3337 24172 3358 24212
rect 3358 24172 3398 24212
rect 3398 24172 3423 24212
rect 3169 24149 3255 24172
rect 3337 24149 3423 24172
rect 18289 24212 18375 24235
rect 18457 24212 18543 24235
rect 18289 24172 18314 24212
rect 18314 24172 18354 24212
rect 18354 24172 18375 24212
rect 18457 24172 18478 24212
rect 18478 24172 18518 24212
rect 18518 24172 18543 24212
rect 18289 24149 18375 24172
rect 18457 24149 18543 24172
rect 33409 24212 33495 24235
rect 33577 24212 33663 24235
rect 33409 24172 33434 24212
rect 33434 24172 33474 24212
rect 33474 24172 33495 24212
rect 33577 24172 33598 24212
rect 33598 24172 33638 24212
rect 33638 24172 33663 24212
rect 33409 24149 33495 24172
rect 33577 24149 33663 24172
rect 48529 24212 48615 24235
rect 48697 24212 48783 24235
rect 48529 24172 48554 24212
rect 48554 24172 48594 24212
rect 48594 24172 48615 24212
rect 48697 24172 48718 24212
rect 48718 24172 48758 24212
rect 48758 24172 48783 24212
rect 48529 24149 48615 24172
rect 48697 24149 48783 24172
rect 63649 24212 63735 24235
rect 63817 24212 63903 24235
rect 63649 24172 63674 24212
rect 63674 24172 63714 24212
rect 63714 24172 63735 24212
rect 63817 24172 63838 24212
rect 63838 24172 63878 24212
rect 63878 24172 63903 24212
rect 63649 24149 63735 24172
rect 63817 24149 63903 24172
rect 78769 24212 78855 24235
rect 78937 24212 79023 24235
rect 78769 24172 78794 24212
rect 78794 24172 78834 24212
rect 78834 24172 78855 24212
rect 78937 24172 78958 24212
rect 78958 24172 78998 24212
rect 78998 24172 79023 24212
rect 78769 24149 78855 24172
rect 78937 24149 79023 24172
rect 93889 24212 93975 24235
rect 94057 24212 94143 24235
rect 93889 24172 93914 24212
rect 93914 24172 93954 24212
rect 93954 24172 93975 24212
rect 94057 24172 94078 24212
rect 94078 24172 94118 24212
rect 94118 24172 94143 24212
rect 93889 24149 93975 24172
rect 94057 24149 94143 24172
rect 4409 23456 4495 23479
rect 4577 23456 4663 23479
rect 4409 23416 4434 23456
rect 4434 23416 4474 23456
rect 4474 23416 4495 23456
rect 4577 23416 4598 23456
rect 4598 23416 4638 23456
rect 4638 23416 4663 23456
rect 4409 23393 4495 23416
rect 4577 23393 4663 23416
rect 19529 23456 19615 23479
rect 19697 23456 19783 23479
rect 19529 23416 19554 23456
rect 19554 23416 19594 23456
rect 19594 23416 19615 23456
rect 19697 23416 19718 23456
rect 19718 23416 19758 23456
rect 19758 23416 19783 23456
rect 19529 23393 19615 23416
rect 19697 23393 19783 23416
rect 34649 23456 34735 23479
rect 34817 23456 34903 23479
rect 34649 23416 34674 23456
rect 34674 23416 34714 23456
rect 34714 23416 34735 23456
rect 34817 23416 34838 23456
rect 34838 23416 34878 23456
rect 34878 23416 34903 23456
rect 34649 23393 34735 23416
rect 34817 23393 34903 23416
rect 49769 23456 49855 23479
rect 49937 23456 50023 23479
rect 49769 23416 49794 23456
rect 49794 23416 49834 23456
rect 49834 23416 49855 23456
rect 49937 23416 49958 23456
rect 49958 23416 49998 23456
rect 49998 23416 50023 23456
rect 49769 23393 49855 23416
rect 49937 23393 50023 23416
rect 64889 23456 64975 23479
rect 65057 23456 65143 23479
rect 64889 23416 64914 23456
rect 64914 23416 64954 23456
rect 64954 23416 64975 23456
rect 65057 23416 65078 23456
rect 65078 23416 65118 23456
rect 65118 23416 65143 23456
rect 64889 23393 64975 23416
rect 65057 23393 65143 23416
rect 80009 23456 80095 23479
rect 80177 23456 80263 23479
rect 80009 23416 80034 23456
rect 80034 23416 80074 23456
rect 80074 23416 80095 23456
rect 80177 23416 80198 23456
rect 80198 23416 80238 23456
rect 80238 23416 80263 23456
rect 80009 23393 80095 23416
rect 80177 23393 80263 23416
rect 95129 23456 95215 23479
rect 95297 23456 95383 23479
rect 95129 23416 95154 23456
rect 95154 23416 95194 23456
rect 95194 23416 95215 23456
rect 95297 23416 95318 23456
rect 95318 23416 95358 23456
rect 95358 23416 95383 23456
rect 95129 23393 95215 23416
rect 95297 23393 95383 23416
rect 3169 22700 3255 22723
rect 3337 22700 3423 22723
rect 3169 22660 3194 22700
rect 3194 22660 3234 22700
rect 3234 22660 3255 22700
rect 3337 22660 3358 22700
rect 3358 22660 3398 22700
rect 3398 22660 3423 22700
rect 3169 22637 3255 22660
rect 3337 22637 3423 22660
rect 18289 22700 18375 22723
rect 18457 22700 18543 22723
rect 18289 22660 18314 22700
rect 18314 22660 18354 22700
rect 18354 22660 18375 22700
rect 18457 22660 18478 22700
rect 18478 22660 18518 22700
rect 18518 22660 18543 22700
rect 18289 22637 18375 22660
rect 18457 22637 18543 22660
rect 33409 22700 33495 22723
rect 33577 22700 33663 22723
rect 33409 22660 33434 22700
rect 33434 22660 33474 22700
rect 33474 22660 33495 22700
rect 33577 22660 33598 22700
rect 33598 22660 33638 22700
rect 33638 22660 33663 22700
rect 33409 22637 33495 22660
rect 33577 22637 33663 22660
rect 48529 22700 48615 22723
rect 48697 22700 48783 22723
rect 48529 22660 48554 22700
rect 48554 22660 48594 22700
rect 48594 22660 48615 22700
rect 48697 22660 48718 22700
rect 48718 22660 48758 22700
rect 48758 22660 48783 22700
rect 48529 22637 48615 22660
rect 48697 22637 48783 22660
rect 63649 22700 63735 22723
rect 63817 22700 63903 22723
rect 63649 22660 63674 22700
rect 63674 22660 63714 22700
rect 63714 22660 63735 22700
rect 63817 22660 63838 22700
rect 63838 22660 63878 22700
rect 63878 22660 63903 22700
rect 63649 22637 63735 22660
rect 63817 22637 63903 22660
rect 78769 22700 78855 22723
rect 78937 22700 79023 22723
rect 78769 22660 78794 22700
rect 78794 22660 78834 22700
rect 78834 22660 78855 22700
rect 78937 22660 78958 22700
rect 78958 22660 78998 22700
rect 78998 22660 79023 22700
rect 78769 22637 78855 22660
rect 78937 22637 79023 22660
rect 93889 22700 93975 22723
rect 94057 22700 94143 22723
rect 93889 22660 93914 22700
rect 93914 22660 93954 22700
rect 93954 22660 93975 22700
rect 94057 22660 94078 22700
rect 94078 22660 94118 22700
rect 94118 22660 94143 22700
rect 93889 22637 93975 22660
rect 94057 22637 94143 22660
rect 4409 21944 4495 21967
rect 4577 21944 4663 21967
rect 4409 21904 4434 21944
rect 4434 21904 4474 21944
rect 4474 21904 4495 21944
rect 4577 21904 4598 21944
rect 4598 21904 4638 21944
rect 4638 21904 4663 21944
rect 4409 21881 4495 21904
rect 4577 21881 4663 21904
rect 19529 21944 19615 21967
rect 19697 21944 19783 21967
rect 19529 21904 19554 21944
rect 19554 21904 19594 21944
rect 19594 21904 19615 21944
rect 19697 21904 19718 21944
rect 19718 21904 19758 21944
rect 19758 21904 19783 21944
rect 19529 21881 19615 21904
rect 19697 21881 19783 21904
rect 34649 21944 34735 21967
rect 34817 21944 34903 21967
rect 34649 21904 34674 21944
rect 34674 21904 34714 21944
rect 34714 21904 34735 21944
rect 34817 21904 34838 21944
rect 34838 21904 34878 21944
rect 34878 21904 34903 21944
rect 34649 21881 34735 21904
rect 34817 21881 34903 21904
rect 49769 21944 49855 21967
rect 49937 21944 50023 21967
rect 49769 21904 49794 21944
rect 49794 21904 49834 21944
rect 49834 21904 49855 21944
rect 49937 21904 49958 21944
rect 49958 21904 49998 21944
rect 49998 21904 50023 21944
rect 49769 21881 49855 21904
rect 49937 21881 50023 21904
rect 64889 21944 64975 21967
rect 65057 21944 65143 21967
rect 64889 21904 64914 21944
rect 64914 21904 64954 21944
rect 64954 21904 64975 21944
rect 65057 21904 65078 21944
rect 65078 21904 65118 21944
rect 65118 21904 65143 21944
rect 64889 21881 64975 21904
rect 65057 21881 65143 21904
rect 80009 21944 80095 21967
rect 80177 21944 80263 21967
rect 80009 21904 80034 21944
rect 80034 21904 80074 21944
rect 80074 21904 80095 21944
rect 80177 21904 80198 21944
rect 80198 21904 80238 21944
rect 80238 21904 80263 21944
rect 80009 21881 80095 21904
rect 80177 21881 80263 21904
rect 95129 21944 95215 21967
rect 95297 21944 95383 21967
rect 95129 21904 95154 21944
rect 95154 21904 95194 21944
rect 95194 21904 95215 21944
rect 95297 21904 95318 21944
rect 95318 21904 95358 21944
rect 95358 21904 95383 21944
rect 95129 21881 95215 21904
rect 95297 21881 95383 21904
rect 3169 21188 3255 21211
rect 3337 21188 3423 21211
rect 3169 21148 3194 21188
rect 3194 21148 3234 21188
rect 3234 21148 3255 21188
rect 3337 21148 3358 21188
rect 3358 21148 3398 21188
rect 3398 21148 3423 21188
rect 3169 21125 3255 21148
rect 3337 21125 3423 21148
rect 18289 21188 18375 21211
rect 18457 21188 18543 21211
rect 18289 21148 18314 21188
rect 18314 21148 18354 21188
rect 18354 21148 18375 21188
rect 18457 21148 18478 21188
rect 18478 21148 18518 21188
rect 18518 21148 18543 21188
rect 18289 21125 18375 21148
rect 18457 21125 18543 21148
rect 33409 21188 33495 21211
rect 33577 21188 33663 21211
rect 33409 21148 33434 21188
rect 33434 21148 33474 21188
rect 33474 21148 33495 21188
rect 33577 21148 33598 21188
rect 33598 21148 33638 21188
rect 33638 21148 33663 21188
rect 33409 21125 33495 21148
rect 33577 21125 33663 21148
rect 48529 21188 48615 21211
rect 48697 21188 48783 21211
rect 48529 21148 48554 21188
rect 48554 21148 48594 21188
rect 48594 21148 48615 21188
rect 48697 21148 48718 21188
rect 48718 21148 48758 21188
rect 48758 21148 48783 21188
rect 48529 21125 48615 21148
rect 48697 21125 48783 21148
rect 63649 21188 63735 21211
rect 63817 21188 63903 21211
rect 63649 21148 63674 21188
rect 63674 21148 63714 21188
rect 63714 21148 63735 21188
rect 63817 21148 63838 21188
rect 63838 21148 63878 21188
rect 63878 21148 63903 21188
rect 63649 21125 63735 21148
rect 63817 21125 63903 21148
rect 78769 21188 78855 21211
rect 78937 21188 79023 21211
rect 78769 21148 78794 21188
rect 78794 21148 78834 21188
rect 78834 21148 78855 21188
rect 78937 21148 78958 21188
rect 78958 21148 78998 21188
rect 78998 21148 79023 21188
rect 78769 21125 78855 21148
rect 78937 21125 79023 21148
rect 93889 21188 93975 21211
rect 94057 21188 94143 21211
rect 93889 21148 93914 21188
rect 93914 21148 93954 21188
rect 93954 21148 93975 21188
rect 94057 21148 94078 21188
rect 94078 21148 94118 21188
rect 94118 21148 94143 21188
rect 93889 21125 93975 21148
rect 94057 21125 94143 21148
rect 4409 20432 4495 20455
rect 4577 20432 4663 20455
rect 4409 20392 4434 20432
rect 4434 20392 4474 20432
rect 4474 20392 4495 20432
rect 4577 20392 4598 20432
rect 4598 20392 4638 20432
rect 4638 20392 4663 20432
rect 4409 20369 4495 20392
rect 4577 20369 4663 20392
rect 19529 20432 19615 20455
rect 19697 20432 19783 20455
rect 19529 20392 19554 20432
rect 19554 20392 19594 20432
rect 19594 20392 19615 20432
rect 19697 20392 19718 20432
rect 19718 20392 19758 20432
rect 19758 20392 19783 20432
rect 19529 20369 19615 20392
rect 19697 20369 19783 20392
rect 34649 20432 34735 20455
rect 34817 20432 34903 20455
rect 34649 20392 34674 20432
rect 34674 20392 34714 20432
rect 34714 20392 34735 20432
rect 34817 20392 34838 20432
rect 34838 20392 34878 20432
rect 34878 20392 34903 20432
rect 34649 20369 34735 20392
rect 34817 20369 34903 20392
rect 49769 20432 49855 20455
rect 49937 20432 50023 20455
rect 49769 20392 49794 20432
rect 49794 20392 49834 20432
rect 49834 20392 49855 20432
rect 49937 20392 49958 20432
rect 49958 20392 49998 20432
rect 49998 20392 50023 20432
rect 49769 20369 49855 20392
rect 49937 20369 50023 20392
rect 64889 20432 64975 20455
rect 65057 20432 65143 20455
rect 64889 20392 64914 20432
rect 64914 20392 64954 20432
rect 64954 20392 64975 20432
rect 65057 20392 65078 20432
rect 65078 20392 65118 20432
rect 65118 20392 65143 20432
rect 64889 20369 64975 20392
rect 65057 20369 65143 20392
rect 80009 20432 80095 20455
rect 80177 20432 80263 20455
rect 80009 20392 80034 20432
rect 80034 20392 80074 20432
rect 80074 20392 80095 20432
rect 80177 20392 80198 20432
rect 80198 20392 80238 20432
rect 80238 20392 80263 20432
rect 80009 20369 80095 20392
rect 80177 20369 80263 20392
rect 95129 20432 95215 20455
rect 95297 20432 95383 20455
rect 95129 20392 95154 20432
rect 95154 20392 95194 20432
rect 95194 20392 95215 20432
rect 95297 20392 95318 20432
rect 95318 20392 95358 20432
rect 95358 20392 95383 20432
rect 95129 20369 95215 20392
rect 95297 20369 95383 20392
rect 3169 19676 3255 19699
rect 3337 19676 3423 19699
rect 3169 19636 3194 19676
rect 3194 19636 3234 19676
rect 3234 19636 3255 19676
rect 3337 19636 3358 19676
rect 3358 19636 3398 19676
rect 3398 19636 3423 19676
rect 3169 19613 3255 19636
rect 3337 19613 3423 19636
rect 18289 19676 18375 19699
rect 18457 19676 18543 19699
rect 18289 19636 18314 19676
rect 18314 19636 18354 19676
rect 18354 19636 18375 19676
rect 18457 19636 18478 19676
rect 18478 19636 18518 19676
rect 18518 19636 18543 19676
rect 18289 19613 18375 19636
rect 18457 19613 18543 19636
rect 33409 19676 33495 19699
rect 33577 19676 33663 19699
rect 33409 19636 33434 19676
rect 33434 19636 33474 19676
rect 33474 19636 33495 19676
rect 33577 19636 33598 19676
rect 33598 19636 33638 19676
rect 33638 19636 33663 19676
rect 33409 19613 33495 19636
rect 33577 19613 33663 19636
rect 48529 19676 48615 19699
rect 48697 19676 48783 19699
rect 48529 19636 48554 19676
rect 48554 19636 48594 19676
rect 48594 19636 48615 19676
rect 48697 19636 48718 19676
rect 48718 19636 48758 19676
rect 48758 19636 48783 19676
rect 48529 19613 48615 19636
rect 48697 19613 48783 19636
rect 63649 19676 63735 19699
rect 63817 19676 63903 19699
rect 63649 19636 63674 19676
rect 63674 19636 63714 19676
rect 63714 19636 63735 19676
rect 63817 19636 63838 19676
rect 63838 19636 63878 19676
rect 63878 19636 63903 19676
rect 63649 19613 63735 19636
rect 63817 19613 63903 19636
rect 78769 19676 78855 19699
rect 78937 19676 79023 19699
rect 78769 19636 78794 19676
rect 78794 19636 78834 19676
rect 78834 19636 78855 19676
rect 78937 19636 78958 19676
rect 78958 19636 78998 19676
rect 78998 19636 79023 19676
rect 78769 19613 78855 19636
rect 78937 19613 79023 19636
rect 93889 19676 93975 19699
rect 94057 19676 94143 19699
rect 93889 19636 93914 19676
rect 93914 19636 93954 19676
rect 93954 19636 93975 19676
rect 94057 19636 94078 19676
rect 94078 19636 94118 19676
rect 94118 19636 94143 19676
rect 93889 19613 93975 19636
rect 94057 19613 94143 19636
rect 4409 18920 4495 18943
rect 4577 18920 4663 18943
rect 4409 18880 4434 18920
rect 4434 18880 4474 18920
rect 4474 18880 4495 18920
rect 4577 18880 4598 18920
rect 4598 18880 4638 18920
rect 4638 18880 4663 18920
rect 4409 18857 4495 18880
rect 4577 18857 4663 18880
rect 19529 18920 19615 18943
rect 19697 18920 19783 18943
rect 19529 18880 19554 18920
rect 19554 18880 19594 18920
rect 19594 18880 19615 18920
rect 19697 18880 19718 18920
rect 19718 18880 19758 18920
rect 19758 18880 19783 18920
rect 19529 18857 19615 18880
rect 19697 18857 19783 18880
rect 34649 18920 34735 18943
rect 34817 18920 34903 18943
rect 34649 18880 34674 18920
rect 34674 18880 34714 18920
rect 34714 18880 34735 18920
rect 34817 18880 34838 18920
rect 34838 18880 34878 18920
rect 34878 18880 34903 18920
rect 34649 18857 34735 18880
rect 34817 18857 34903 18880
rect 49769 18920 49855 18943
rect 49937 18920 50023 18943
rect 49769 18880 49794 18920
rect 49794 18880 49834 18920
rect 49834 18880 49855 18920
rect 49937 18880 49958 18920
rect 49958 18880 49998 18920
rect 49998 18880 50023 18920
rect 49769 18857 49855 18880
rect 49937 18857 50023 18880
rect 64889 18920 64975 18943
rect 65057 18920 65143 18943
rect 64889 18880 64914 18920
rect 64914 18880 64954 18920
rect 64954 18880 64975 18920
rect 65057 18880 65078 18920
rect 65078 18880 65118 18920
rect 65118 18880 65143 18920
rect 64889 18857 64975 18880
rect 65057 18857 65143 18880
rect 80009 18920 80095 18943
rect 80177 18920 80263 18943
rect 80009 18880 80034 18920
rect 80034 18880 80074 18920
rect 80074 18880 80095 18920
rect 80177 18880 80198 18920
rect 80198 18880 80238 18920
rect 80238 18880 80263 18920
rect 80009 18857 80095 18880
rect 80177 18857 80263 18880
rect 95129 18920 95215 18943
rect 95297 18920 95383 18943
rect 95129 18880 95154 18920
rect 95154 18880 95194 18920
rect 95194 18880 95215 18920
rect 95297 18880 95318 18920
rect 95318 18880 95358 18920
rect 95358 18880 95383 18920
rect 95129 18857 95215 18880
rect 95297 18857 95383 18880
rect 3169 18164 3255 18187
rect 3337 18164 3423 18187
rect 3169 18124 3194 18164
rect 3194 18124 3234 18164
rect 3234 18124 3255 18164
rect 3337 18124 3358 18164
rect 3358 18124 3398 18164
rect 3398 18124 3423 18164
rect 3169 18101 3255 18124
rect 3337 18101 3423 18124
rect 18289 18164 18375 18187
rect 18457 18164 18543 18187
rect 18289 18124 18314 18164
rect 18314 18124 18354 18164
rect 18354 18124 18375 18164
rect 18457 18124 18478 18164
rect 18478 18124 18518 18164
rect 18518 18124 18543 18164
rect 18289 18101 18375 18124
rect 18457 18101 18543 18124
rect 33409 18164 33495 18187
rect 33577 18164 33663 18187
rect 33409 18124 33434 18164
rect 33434 18124 33474 18164
rect 33474 18124 33495 18164
rect 33577 18124 33598 18164
rect 33598 18124 33638 18164
rect 33638 18124 33663 18164
rect 33409 18101 33495 18124
rect 33577 18101 33663 18124
rect 48529 18164 48615 18187
rect 48697 18164 48783 18187
rect 48529 18124 48554 18164
rect 48554 18124 48594 18164
rect 48594 18124 48615 18164
rect 48697 18124 48718 18164
rect 48718 18124 48758 18164
rect 48758 18124 48783 18164
rect 48529 18101 48615 18124
rect 48697 18101 48783 18124
rect 63649 18164 63735 18187
rect 63817 18164 63903 18187
rect 63649 18124 63674 18164
rect 63674 18124 63714 18164
rect 63714 18124 63735 18164
rect 63817 18124 63838 18164
rect 63838 18124 63878 18164
rect 63878 18124 63903 18164
rect 63649 18101 63735 18124
rect 63817 18101 63903 18124
rect 78769 18164 78855 18187
rect 78937 18164 79023 18187
rect 78769 18124 78794 18164
rect 78794 18124 78834 18164
rect 78834 18124 78855 18164
rect 78937 18124 78958 18164
rect 78958 18124 78998 18164
rect 78998 18124 79023 18164
rect 78769 18101 78855 18124
rect 78937 18101 79023 18124
rect 93889 18164 93975 18187
rect 94057 18164 94143 18187
rect 93889 18124 93914 18164
rect 93914 18124 93954 18164
rect 93954 18124 93975 18164
rect 94057 18124 94078 18164
rect 94078 18124 94118 18164
rect 94118 18124 94143 18164
rect 93889 18101 93975 18124
rect 94057 18101 94143 18124
rect 4409 17408 4495 17431
rect 4577 17408 4663 17431
rect 4409 17368 4434 17408
rect 4434 17368 4474 17408
rect 4474 17368 4495 17408
rect 4577 17368 4598 17408
rect 4598 17368 4638 17408
rect 4638 17368 4663 17408
rect 4409 17345 4495 17368
rect 4577 17345 4663 17368
rect 19529 17408 19615 17431
rect 19697 17408 19783 17431
rect 19529 17368 19554 17408
rect 19554 17368 19594 17408
rect 19594 17368 19615 17408
rect 19697 17368 19718 17408
rect 19718 17368 19758 17408
rect 19758 17368 19783 17408
rect 19529 17345 19615 17368
rect 19697 17345 19783 17368
rect 34649 17408 34735 17431
rect 34817 17408 34903 17431
rect 34649 17368 34674 17408
rect 34674 17368 34714 17408
rect 34714 17368 34735 17408
rect 34817 17368 34838 17408
rect 34838 17368 34878 17408
rect 34878 17368 34903 17408
rect 34649 17345 34735 17368
rect 34817 17345 34903 17368
rect 49769 17408 49855 17431
rect 49937 17408 50023 17431
rect 49769 17368 49794 17408
rect 49794 17368 49834 17408
rect 49834 17368 49855 17408
rect 49937 17368 49958 17408
rect 49958 17368 49998 17408
rect 49998 17368 50023 17408
rect 49769 17345 49855 17368
rect 49937 17345 50023 17368
rect 64889 17408 64975 17431
rect 65057 17408 65143 17431
rect 64889 17368 64914 17408
rect 64914 17368 64954 17408
rect 64954 17368 64975 17408
rect 65057 17368 65078 17408
rect 65078 17368 65118 17408
rect 65118 17368 65143 17408
rect 64889 17345 64975 17368
rect 65057 17345 65143 17368
rect 80009 17408 80095 17431
rect 80177 17408 80263 17431
rect 80009 17368 80034 17408
rect 80034 17368 80074 17408
rect 80074 17368 80095 17408
rect 80177 17368 80198 17408
rect 80198 17368 80238 17408
rect 80238 17368 80263 17408
rect 80009 17345 80095 17368
rect 80177 17345 80263 17368
rect 95129 17408 95215 17431
rect 95297 17408 95383 17431
rect 95129 17368 95154 17408
rect 95154 17368 95194 17408
rect 95194 17368 95215 17408
rect 95297 17368 95318 17408
rect 95318 17368 95358 17408
rect 95358 17368 95383 17408
rect 95129 17345 95215 17368
rect 95297 17345 95383 17368
rect 3169 16652 3255 16675
rect 3337 16652 3423 16675
rect 3169 16612 3194 16652
rect 3194 16612 3234 16652
rect 3234 16612 3255 16652
rect 3337 16612 3358 16652
rect 3358 16612 3398 16652
rect 3398 16612 3423 16652
rect 3169 16589 3255 16612
rect 3337 16589 3423 16612
rect 18289 16652 18375 16675
rect 18457 16652 18543 16675
rect 18289 16612 18314 16652
rect 18314 16612 18354 16652
rect 18354 16612 18375 16652
rect 18457 16612 18478 16652
rect 18478 16612 18518 16652
rect 18518 16612 18543 16652
rect 18289 16589 18375 16612
rect 18457 16589 18543 16612
rect 33409 16652 33495 16675
rect 33577 16652 33663 16675
rect 33409 16612 33434 16652
rect 33434 16612 33474 16652
rect 33474 16612 33495 16652
rect 33577 16612 33598 16652
rect 33598 16612 33638 16652
rect 33638 16612 33663 16652
rect 33409 16589 33495 16612
rect 33577 16589 33663 16612
rect 48529 16652 48615 16675
rect 48697 16652 48783 16675
rect 48529 16612 48554 16652
rect 48554 16612 48594 16652
rect 48594 16612 48615 16652
rect 48697 16612 48718 16652
rect 48718 16612 48758 16652
rect 48758 16612 48783 16652
rect 48529 16589 48615 16612
rect 48697 16589 48783 16612
rect 63649 16652 63735 16675
rect 63817 16652 63903 16675
rect 63649 16612 63674 16652
rect 63674 16612 63714 16652
rect 63714 16612 63735 16652
rect 63817 16612 63838 16652
rect 63838 16612 63878 16652
rect 63878 16612 63903 16652
rect 63649 16589 63735 16612
rect 63817 16589 63903 16612
rect 78769 16652 78855 16675
rect 78937 16652 79023 16675
rect 78769 16612 78794 16652
rect 78794 16612 78834 16652
rect 78834 16612 78855 16652
rect 78937 16612 78958 16652
rect 78958 16612 78998 16652
rect 78998 16612 79023 16652
rect 78769 16589 78855 16612
rect 78937 16589 79023 16612
rect 93889 16652 93975 16675
rect 94057 16652 94143 16675
rect 93889 16612 93914 16652
rect 93914 16612 93954 16652
rect 93954 16612 93975 16652
rect 94057 16612 94078 16652
rect 94078 16612 94118 16652
rect 94118 16612 94143 16652
rect 93889 16589 93975 16612
rect 94057 16589 94143 16612
rect 4409 15896 4495 15919
rect 4577 15896 4663 15919
rect 4409 15856 4434 15896
rect 4434 15856 4474 15896
rect 4474 15856 4495 15896
rect 4577 15856 4598 15896
rect 4598 15856 4638 15896
rect 4638 15856 4663 15896
rect 4409 15833 4495 15856
rect 4577 15833 4663 15856
rect 19529 15896 19615 15919
rect 19697 15896 19783 15919
rect 19529 15856 19554 15896
rect 19554 15856 19594 15896
rect 19594 15856 19615 15896
rect 19697 15856 19718 15896
rect 19718 15856 19758 15896
rect 19758 15856 19783 15896
rect 19529 15833 19615 15856
rect 19697 15833 19783 15856
rect 34649 15896 34735 15919
rect 34817 15896 34903 15919
rect 34649 15856 34674 15896
rect 34674 15856 34714 15896
rect 34714 15856 34735 15896
rect 34817 15856 34838 15896
rect 34838 15856 34878 15896
rect 34878 15856 34903 15896
rect 34649 15833 34735 15856
rect 34817 15833 34903 15856
rect 49769 15896 49855 15919
rect 49937 15896 50023 15919
rect 49769 15856 49794 15896
rect 49794 15856 49834 15896
rect 49834 15856 49855 15896
rect 49937 15856 49958 15896
rect 49958 15856 49998 15896
rect 49998 15856 50023 15896
rect 49769 15833 49855 15856
rect 49937 15833 50023 15856
rect 64889 15896 64975 15919
rect 65057 15896 65143 15919
rect 64889 15856 64914 15896
rect 64914 15856 64954 15896
rect 64954 15856 64975 15896
rect 65057 15856 65078 15896
rect 65078 15856 65118 15896
rect 65118 15856 65143 15896
rect 64889 15833 64975 15856
rect 65057 15833 65143 15856
rect 80009 15896 80095 15919
rect 80177 15896 80263 15919
rect 80009 15856 80034 15896
rect 80034 15856 80074 15896
rect 80074 15856 80095 15896
rect 80177 15856 80198 15896
rect 80198 15856 80238 15896
rect 80238 15856 80263 15896
rect 80009 15833 80095 15856
rect 80177 15833 80263 15856
rect 95129 15896 95215 15919
rect 95297 15896 95383 15919
rect 95129 15856 95154 15896
rect 95154 15856 95194 15896
rect 95194 15856 95215 15896
rect 95297 15856 95318 15896
rect 95318 15856 95358 15896
rect 95358 15856 95383 15896
rect 95129 15833 95215 15856
rect 95297 15833 95383 15856
rect 3169 15140 3255 15163
rect 3337 15140 3423 15163
rect 3169 15100 3194 15140
rect 3194 15100 3234 15140
rect 3234 15100 3255 15140
rect 3337 15100 3358 15140
rect 3358 15100 3398 15140
rect 3398 15100 3423 15140
rect 3169 15077 3255 15100
rect 3337 15077 3423 15100
rect 18289 15140 18375 15163
rect 18457 15140 18543 15163
rect 18289 15100 18314 15140
rect 18314 15100 18354 15140
rect 18354 15100 18375 15140
rect 18457 15100 18478 15140
rect 18478 15100 18518 15140
rect 18518 15100 18543 15140
rect 18289 15077 18375 15100
rect 18457 15077 18543 15100
rect 33409 15140 33495 15163
rect 33577 15140 33663 15163
rect 33409 15100 33434 15140
rect 33434 15100 33474 15140
rect 33474 15100 33495 15140
rect 33577 15100 33598 15140
rect 33598 15100 33638 15140
rect 33638 15100 33663 15140
rect 33409 15077 33495 15100
rect 33577 15077 33663 15100
rect 48529 15140 48615 15163
rect 48697 15140 48783 15163
rect 48529 15100 48554 15140
rect 48554 15100 48594 15140
rect 48594 15100 48615 15140
rect 48697 15100 48718 15140
rect 48718 15100 48758 15140
rect 48758 15100 48783 15140
rect 48529 15077 48615 15100
rect 48697 15077 48783 15100
rect 63649 15140 63735 15163
rect 63817 15140 63903 15163
rect 63649 15100 63674 15140
rect 63674 15100 63714 15140
rect 63714 15100 63735 15140
rect 63817 15100 63838 15140
rect 63838 15100 63878 15140
rect 63878 15100 63903 15140
rect 63649 15077 63735 15100
rect 63817 15077 63903 15100
rect 78769 15140 78855 15163
rect 78937 15140 79023 15163
rect 78769 15100 78794 15140
rect 78794 15100 78834 15140
rect 78834 15100 78855 15140
rect 78937 15100 78958 15140
rect 78958 15100 78998 15140
rect 78998 15100 79023 15140
rect 78769 15077 78855 15100
rect 78937 15077 79023 15100
rect 93889 15140 93975 15163
rect 94057 15140 94143 15163
rect 93889 15100 93914 15140
rect 93914 15100 93954 15140
rect 93954 15100 93975 15140
rect 94057 15100 94078 15140
rect 94078 15100 94118 15140
rect 94118 15100 94143 15140
rect 93889 15077 93975 15100
rect 94057 15077 94143 15100
rect 4409 14384 4495 14407
rect 4577 14384 4663 14407
rect 4409 14344 4434 14384
rect 4434 14344 4474 14384
rect 4474 14344 4495 14384
rect 4577 14344 4598 14384
rect 4598 14344 4638 14384
rect 4638 14344 4663 14384
rect 4409 14321 4495 14344
rect 4577 14321 4663 14344
rect 19529 14384 19615 14407
rect 19697 14384 19783 14407
rect 19529 14344 19554 14384
rect 19554 14344 19594 14384
rect 19594 14344 19615 14384
rect 19697 14344 19718 14384
rect 19718 14344 19758 14384
rect 19758 14344 19783 14384
rect 19529 14321 19615 14344
rect 19697 14321 19783 14344
rect 34649 14384 34735 14407
rect 34817 14384 34903 14407
rect 34649 14344 34674 14384
rect 34674 14344 34714 14384
rect 34714 14344 34735 14384
rect 34817 14344 34838 14384
rect 34838 14344 34878 14384
rect 34878 14344 34903 14384
rect 34649 14321 34735 14344
rect 34817 14321 34903 14344
rect 49769 14384 49855 14407
rect 49937 14384 50023 14407
rect 49769 14344 49794 14384
rect 49794 14344 49834 14384
rect 49834 14344 49855 14384
rect 49937 14344 49958 14384
rect 49958 14344 49998 14384
rect 49998 14344 50023 14384
rect 49769 14321 49855 14344
rect 49937 14321 50023 14344
rect 64889 14384 64975 14407
rect 65057 14384 65143 14407
rect 64889 14344 64914 14384
rect 64914 14344 64954 14384
rect 64954 14344 64975 14384
rect 65057 14344 65078 14384
rect 65078 14344 65118 14384
rect 65118 14344 65143 14384
rect 64889 14321 64975 14344
rect 65057 14321 65143 14344
rect 80009 14384 80095 14407
rect 80177 14384 80263 14407
rect 80009 14344 80034 14384
rect 80034 14344 80074 14384
rect 80074 14344 80095 14384
rect 80177 14344 80198 14384
rect 80198 14344 80238 14384
rect 80238 14344 80263 14384
rect 80009 14321 80095 14344
rect 80177 14321 80263 14344
rect 95129 14384 95215 14407
rect 95297 14384 95383 14407
rect 95129 14344 95154 14384
rect 95154 14344 95194 14384
rect 95194 14344 95215 14384
rect 95297 14344 95318 14384
rect 95318 14344 95358 14384
rect 95358 14344 95383 14384
rect 95129 14321 95215 14344
rect 95297 14321 95383 14344
rect 3169 13628 3255 13651
rect 3337 13628 3423 13651
rect 3169 13588 3194 13628
rect 3194 13588 3234 13628
rect 3234 13588 3255 13628
rect 3337 13588 3358 13628
rect 3358 13588 3398 13628
rect 3398 13588 3423 13628
rect 3169 13565 3255 13588
rect 3337 13565 3423 13588
rect 18289 13628 18375 13651
rect 18457 13628 18543 13651
rect 18289 13588 18314 13628
rect 18314 13588 18354 13628
rect 18354 13588 18375 13628
rect 18457 13588 18478 13628
rect 18478 13588 18518 13628
rect 18518 13588 18543 13628
rect 18289 13565 18375 13588
rect 18457 13565 18543 13588
rect 33409 13628 33495 13651
rect 33577 13628 33663 13651
rect 33409 13588 33434 13628
rect 33434 13588 33474 13628
rect 33474 13588 33495 13628
rect 33577 13588 33598 13628
rect 33598 13588 33638 13628
rect 33638 13588 33663 13628
rect 33409 13565 33495 13588
rect 33577 13565 33663 13588
rect 48529 13628 48615 13651
rect 48697 13628 48783 13651
rect 48529 13588 48554 13628
rect 48554 13588 48594 13628
rect 48594 13588 48615 13628
rect 48697 13588 48718 13628
rect 48718 13588 48758 13628
rect 48758 13588 48783 13628
rect 48529 13565 48615 13588
rect 48697 13565 48783 13588
rect 63649 13628 63735 13651
rect 63817 13628 63903 13651
rect 63649 13588 63674 13628
rect 63674 13588 63714 13628
rect 63714 13588 63735 13628
rect 63817 13588 63838 13628
rect 63838 13588 63878 13628
rect 63878 13588 63903 13628
rect 63649 13565 63735 13588
rect 63817 13565 63903 13588
rect 78769 13628 78855 13651
rect 78937 13628 79023 13651
rect 78769 13588 78794 13628
rect 78794 13588 78834 13628
rect 78834 13588 78855 13628
rect 78937 13588 78958 13628
rect 78958 13588 78998 13628
rect 78998 13588 79023 13628
rect 78769 13565 78855 13588
rect 78937 13565 79023 13588
rect 93889 13628 93975 13651
rect 94057 13628 94143 13651
rect 93889 13588 93914 13628
rect 93914 13588 93954 13628
rect 93954 13588 93975 13628
rect 94057 13588 94078 13628
rect 94078 13588 94118 13628
rect 94118 13588 94143 13628
rect 93889 13565 93975 13588
rect 94057 13565 94143 13588
rect 4409 12872 4495 12895
rect 4577 12872 4663 12895
rect 4409 12832 4434 12872
rect 4434 12832 4474 12872
rect 4474 12832 4495 12872
rect 4577 12832 4598 12872
rect 4598 12832 4638 12872
rect 4638 12832 4663 12872
rect 4409 12809 4495 12832
rect 4577 12809 4663 12832
rect 19529 12872 19615 12895
rect 19697 12872 19783 12895
rect 19529 12832 19554 12872
rect 19554 12832 19594 12872
rect 19594 12832 19615 12872
rect 19697 12832 19718 12872
rect 19718 12832 19758 12872
rect 19758 12832 19783 12872
rect 19529 12809 19615 12832
rect 19697 12809 19783 12832
rect 34649 12872 34735 12895
rect 34817 12872 34903 12895
rect 34649 12832 34674 12872
rect 34674 12832 34714 12872
rect 34714 12832 34735 12872
rect 34817 12832 34838 12872
rect 34838 12832 34878 12872
rect 34878 12832 34903 12872
rect 34649 12809 34735 12832
rect 34817 12809 34903 12832
rect 49769 12872 49855 12895
rect 49937 12872 50023 12895
rect 49769 12832 49794 12872
rect 49794 12832 49834 12872
rect 49834 12832 49855 12872
rect 49937 12832 49958 12872
rect 49958 12832 49998 12872
rect 49998 12832 50023 12872
rect 49769 12809 49855 12832
rect 49937 12809 50023 12832
rect 64889 12872 64975 12895
rect 65057 12872 65143 12895
rect 64889 12832 64914 12872
rect 64914 12832 64954 12872
rect 64954 12832 64975 12872
rect 65057 12832 65078 12872
rect 65078 12832 65118 12872
rect 65118 12832 65143 12872
rect 64889 12809 64975 12832
rect 65057 12809 65143 12832
rect 80009 12872 80095 12895
rect 80177 12872 80263 12895
rect 80009 12832 80034 12872
rect 80034 12832 80074 12872
rect 80074 12832 80095 12872
rect 80177 12832 80198 12872
rect 80198 12832 80238 12872
rect 80238 12832 80263 12872
rect 80009 12809 80095 12832
rect 80177 12809 80263 12832
rect 95129 12872 95215 12895
rect 95297 12872 95383 12895
rect 95129 12832 95154 12872
rect 95154 12832 95194 12872
rect 95194 12832 95215 12872
rect 95297 12832 95318 12872
rect 95318 12832 95358 12872
rect 95358 12832 95383 12872
rect 95129 12809 95215 12832
rect 95297 12809 95383 12832
rect 3169 12116 3255 12139
rect 3337 12116 3423 12139
rect 3169 12076 3194 12116
rect 3194 12076 3234 12116
rect 3234 12076 3255 12116
rect 3337 12076 3358 12116
rect 3358 12076 3398 12116
rect 3398 12076 3423 12116
rect 3169 12053 3255 12076
rect 3337 12053 3423 12076
rect 18289 12116 18375 12139
rect 18457 12116 18543 12139
rect 18289 12076 18314 12116
rect 18314 12076 18354 12116
rect 18354 12076 18375 12116
rect 18457 12076 18478 12116
rect 18478 12076 18518 12116
rect 18518 12076 18543 12116
rect 18289 12053 18375 12076
rect 18457 12053 18543 12076
rect 33409 12116 33495 12139
rect 33577 12116 33663 12139
rect 33409 12076 33434 12116
rect 33434 12076 33474 12116
rect 33474 12076 33495 12116
rect 33577 12076 33598 12116
rect 33598 12076 33638 12116
rect 33638 12076 33663 12116
rect 33409 12053 33495 12076
rect 33577 12053 33663 12076
rect 48529 12116 48615 12139
rect 48697 12116 48783 12139
rect 48529 12076 48554 12116
rect 48554 12076 48594 12116
rect 48594 12076 48615 12116
rect 48697 12076 48718 12116
rect 48718 12076 48758 12116
rect 48758 12076 48783 12116
rect 48529 12053 48615 12076
rect 48697 12053 48783 12076
rect 63649 12116 63735 12139
rect 63817 12116 63903 12139
rect 63649 12076 63674 12116
rect 63674 12076 63714 12116
rect 63714 12076 63735 12116
rect 63817 12076 63838 12116
rect 63838 12076 63878 12116
rect 63878 12076 63903 12116
rect 63649 12053 63735 12076
rect 63817 12053 63903 12076
rect 78769 12116 78855 12139
rect 78937 12116 79023 12139
rect 78769 12076 78794 12116
rect 78794 12076 78834 12116
rect 78834 12076 78855 12116
rect 78937 12076 78958 12116
rect 78958 12076 78998 12116
rect 78998 12076 79023 12116
rect 78769 12053 78855 12076
rect 78937 12053 79023 12076
rect 93889 12116 93975 12139
rect 94057 12116 94143 12139
rect 93889 12076 93914 12116
rect 93914 12076 93954 12116
rect 93954 12076 93975 12116
rect 94057 12076 94078 12116
rect 94078 12076 94118 12116
rect 94118 12076 94143 12116
rect 93889 12053 93975 12076
rect 94057 12053 94143 12076
rect 4409 11360 4495 11383
rect 4577 11360 4663 11383
rect 4409 11320 4434 11360
rect 4434 11320 4474 11360
rect 4474 11320 4495 11360
rect 4577 11320 4598 11360
rect 4598 11320 4638 11360
rect 4638 11320 4663 11360
rect 4409 11297 4495 11320
rect 4577 11297 4663 11320
rect 19529 11360 19615 11383
rect 19697 11360 19783 11383
rect 19529 11320 19554 11360
rect 19554 11320 19594 11360
rect 19594 11320 19615 11360
rect 19697 11320 19718 11360
rect 19718 11320 19758 11360
rect 19758 11320 19783 11360
rect 19529 11297 19615 11320
rect 19697 11297 19783 11320
rect 34649 11360 34735 11383
rect 34817 11360 34903 11383
rect 34649 11320 34674 11360
rect 34674 11320 34714 11360
rect 34714 11320 34735 11360
rect 34817 11320 34838 11360
rect 34838 11320 34878 11360
rect 34878 11320 34903 11360
rect 34649 11297 34735 11320
rect 34817 11297 34903 11320
rect 49769 11360 49855 11383
rect 49937 11360 50023 11383
rect 49769 11320 49794 11360
rect 49794 11320 49834 11360
rect 49834 11320 49855 11360
rect 49937 11320 49958 11360
rect 49958 11320 49998 11360
rect 49998 11320 50023 11360
rect 49769 11297 49855 11320
rect 49937 11297 50023 11320
rect 64889 11360 64975 11383
rect 65057 11360 65143 11383
rect 64889 11320 64914 11360
rect 64914 11320 64954 11360
rect 64954 11320 64975 11360
rect 65057 11320 65078 11360
rect 65078 11320 65118 11360
rect 65118 11320 65143 11360
rect 64889 11297 64975 11320
rect 65057 11297 65143 11320
rect 80009 11360 80095 11383
rect 80177 11360 80263 11383
rect 80009 11320 80034 11360
rect 80034 11320 80074 11360
rect 80074 11320 80095 11360
rect 80177 11320 80198 11360
rect 80198 11320 80238 11360
rect 80238 11320 80263 11360
rect 80009 11297 80095 11320
rect 80177 11297 80263 11320
rect 95129 11360 95215 11383
rect 95297 11360 95383 11383
rect 95129 11320 95154 11360
rect 95154 11320 95194 11360
rect 95194 11320 95215 11360
rect 95297 11320 95318 11360
rect 95318 11320 95358 11360
rect 95358 11320 95383 11360
rect 95129 11297 95215 11320
rect 95297 11297 95383 11320
rect 3169 10604 3255 10627
rect 3337 10604 3423 10627
rect 3169 10564 3194 10604
rect 3194 10564 3234 10604
rect 3234 10564 3255 10604
rect 3337 10564 3358 10604
rect 3358 10564 3398 10604
rect 3398 10564 3423 10604
rect 3169 10541 3255 10564
rect 3337 10541 3423 10564
rect 18289 10604 18375 10627
rect 18457 10604 18543 10627
rect 18289 10564 18314 10604
rect 18314 10564 18354 10604
rect 18354 10564 18375 10604
rect 18457 10564 18478 10604
rect 18478 10564 18518 10604
rect 18518 10564 18543 10604
rect 18289 10541 18375 10564
rect 18457 10541 18543 10564
rect 33409 10604 33495 10627
rect 33577 10604 33663 10627
rect 33409 10564 33434 10604
rect 33434 10564 33474 10604
rect 33474 10564 33495 10604
rect 33577 10564 33598 10604
rect 33598 10564 33638 10604
rect 33638 10564 33663 10604
rect 33409 10541 33495 10564
rect 33577 10541 33663 10564
rect 48529 10604 48615 10627
rect 48697 10604 48783 10627
rect 48529 10564 48554 10604
rect 48554 10564 48594 10604
rect 48594 10564 48615 10604
rect 48697 10564 48718 10604
rect 48718 10564 48758 10604
rect 48758 10564 48783 10604
rect 48529 10541 48615 10564
rect 48697 10541 48783 10564
rect 63649 10604 63735 10627
rect 63817 10604 63903 10627
rect 63649 10564 63674 10604
rect 63674 10564 63714 10604
rect 63714 10564 63735 10604
rect 63817 10564 63838 10604
rect 63838 10564 63878 10604
rect 63878 10564 63903 10604
rect 63649 10541 63735 10564
rect 63817 10541 63903 10564
rect 78769 10604 78855 10627
rect 78937 10604 79023 10627
rect 78769 10564 78794 10604
rect 78794 10564 78834 10604
rect 78834 10564 78855 10604
rect 78937 10564 78958 10604
rect 78958 10564 78998 10604
rect 78998 10564 79023 10604
rect 78769 10541 78855 10564
rect 78937 10541 79023 10564
rect 93889 10604 93975 10627
rect 94057 10604 94143 10627
rect 93889 10564 93914 10604
rect 93914 10564 93954 10604
rect 93954 10564 93975 10604
rect 94057 10564 94078 10604
rect 94078 10564 94118 10604
rect 94118 10564 94143 10604
rect 93889 10541 93975 10564
rect 94057 10541 94143 10564
rect 4409 9848 4495 9871
rect 4577 9848 4663 9871
rect 4409 9808 4434 9848
rect 4434 9808 4474 9848
rect 4474 9808 4495 9848
rect 4577 9808 4598 9848
rect 4598 9808 4638 9848
rect 4638 9808 4663 9848
rect 4409 9785 4495 9808
rect 4577 9785 4663 9808
rect 19529 9848 19615 9871
rect 19697 9848 19783 9871
rect 19529 9808 19554 9848
rect 19554 9808 19594 9848
rect 19594 9808 19615 9848
rect 19697 9808 19718 9848
rect 19718 9808 19758 9848
rect 19758 9808 19783 9848
rect 19529 9785 19615 9808
rect 19697 9785 19783 9808
rect 34649 9848 34735 9871
rect 34817 9848 34903 9871
rect 34649 9808 34674 9848
rect 34674 9808 34714 9848
rect 34714 9808 34735 9848
rect 34817 9808 34838 9848
rect 34838 9808 34878 9848
rect 34878 9808 34903 9848
rect 34649 9785 34735 9808
rect 34817 9785 34903 9808
rect 49769 9848 49855 9871
rect 49937 9848 50023 9871
rect 49769 9808 49794 9848
rect 49794 9808 49834 9848
rect 49834 9808 49855 9848
rect 49937 9808 49958 9848
rect 49958 9808 49998 9848
rect 49998 9808 50023 9848
rect 49769 9785 49855 9808
rect 49937 9785 50023 9808
rect 64889 9848 64975 9871
rect 65057 9848 65143 9871
rect 64889 9808 64914 9848
rect 64914 9808 64954 9848
rect 64954 9808 64975 9848
rect 65057 9808 65078 9848
rect 65078 9808 65118 9848
rect 65118 9808 65143 9848
rect 64889 9785 64975 9808
rect 65057 9785 65143 9808
rect 80009 9848 80095 9871
rect 80177 9848 80263 9871
rect 80009 9808 80034 9848
rect 80034 9808 80074 9848
rect 80074 9808 80095 9848
rect 80177 9808 80198 9848
rect 80198 9808 80238 9848
rect 80238 9808 80263 9848
rect 80009 9785 80095 9808
rect 80177 9785 80263 9808
rect 95129 9848 95215 9871
rect 95297 9848 95383 9871
rect 95129 9808 95154 9848
rect 95154 9808 95194 9848
rect 95194 9808 95215 9848
rect 95297 9808 95318 9848
rect 95318 9808 95358 9848
rect 95358 9808 95383 9848
rect 95129 9785 95215 9808
rect 95297 9785 95383 9808
rect 3169 9092 3255 9115
rect 3337 9092 3423 9115
rect 3169 9052 3194 9092
rect 3194 9052 3234 9092
rect 3234 9052 3255 9092
rect 3337 9052 3358 9092
rect 3358 9052 3398 9092
rect 3398 9052 3423 9092
rect 3169 9029 3255 9052
rect 3337 9029 3423 9052
rect 18289 9092 18375 9115
rect 18457 9092 18543 9115
rect 18289 9052 18314 9092
rect 18314 9052 18354 9092
rect 18354 9052 18375 9092
rect 18457 9052 18478 9092
rect 18478 9052 18518 9092
rect 18518 9052 18543 9092
rect 18289 9029 18375 9052
rect 18457 9029 18543 9052
rect 33409 9092 33495 9115
rect 33577 9092 33663 9115
rect 33409 9052 33434 9092
rect 33434 9052 33474 9092
rect 33474 9052 33495 9092
rect 33577 9052 33598 9092
rect 33598 9052 33638 9092
rect 33638 9052 33663 9092
rect 33409 9029 33495 9052
rect 33577 9029 33663 9052
rect 48529 9092 48615 9115
rect 48697 9092 48783 9115
rect 48529 9052 48554 9092
rect 48554 9052 48594 9092
rect 48594 9052 48615 9092
rect 48697 9052 48718 9092
rect 48718 9052 48758 9092
rect 48758 9052 48783 9092
rect 48529 9029 48615 9052
rect 48697 9029 48783 9052
rect 63649 9092 63735 9115
rect 63817 9092 63903 9115
rect 63649 9052 63674 9092
rect 63674 9052 63714 9092
rect 63714 9052 63735 9092
rect 63817 9052 63838 9092
rect 63838 9052 63878 9092
rect 63878 9052 63903 9092
rect 63649 9029 63735 9052
rect 63817 9029 63903 9052
rect 78769 9092 78855 9115
rect 78937 9092 79023 9115
rect 78769 9052 78794 9092
rect 78794 9052 78834 9092
rect 78834 9052 78855 9092
rect 78937 9052 78958 9092
rect 78958 9052 78998 9092
rect 78998 9052 79023 9092
rect 78769 9029 78855 9052
rect 78937 9029 79023 9052
rect 93889 9092 93975 9115
rect 94057 9092 94143 9115
rect 93889 9052 93914 9092
rect 93914 9052 93954 9092
rect 93954 9052 93975 9092
rect 94057 9052 94078 9092
rect 94078 9052 94118 9092
rect 94118 9052 94143 9092
rect 93889 9029 93975 9052
rect 94057 9029 94143 9052
rect 4409 8336 4495 8359
rect 4577 8336 4663 8359
rect 4409 8296 4434 8336
rect 4434 8296 4474 8336
rect 4474 8296 4495 8336
rect 4577 8296 4598 8336
rect 4598 8296 4638 8336
rect 4638 8296 4663 8336
rect 4409 8273 4495 8296
rect 4577 8273 4663 8296
rect 19529 8336 19615 8359
rect 19697 8336 19783 8359
rect 19529 8296 19554 8336
rect 19554 8296 19594 8336
rect 19594 8296 19615 8336
rect 19697 8296 19718 8336
rect 19718 8296 19758 8336
rect 19758 8296 19783 8336
rect 19529 8273 19615 8296
rect 19697 8273 19783 8296
rect 34649 8336 34735 8359
rect 34817 8336 34903 8359
rect 34649 8296 34674 8336
rect 34674 8296 34714 8336
rect 34714 8296 34735 8336
rect 34817 8296 34838 8336
rect 34838 8296 34878 8336
rect 34878 8296 34903 8336
rect 34649 8273 34735 8296
rect 34817 8273 34903 8296
rect 49769 8336 49855 8359
rect 49937 8336 50023 8359
rect 49769 8296 49794 8336
rect 49794 8296 49834 8336
rect 49834 8296 49855 8336
rect 49937 8296 49958 8336
rect 49958 8296 49998 8336
rect 49998 8296 50023 8336
rect 49769 8273 49855 8296
rect 49937 8273 50023 8296
rect 64889 8336 64975 8359
rect 65057 8336 65143 8359
rect 64889 8296 64914 8336
rect 64914 8296 64954 8336
rect 64954 8296 64975 8336
rect 65057 8296 65078 8336
rect 65078 8296 65118 8336
rect 65118 8296 65143 8336
rect 64889 8273 64975 8296
rect 65057 8273 65143 8296
rect 80009 8336 80095 8359
rect 80177 8336 80263 8359
rect 80009 8296 80034 8336
rect 80034 8296 80074 8336
rect 80074 8296 80095 8336
rect 80177 8296 80198 8336
rect 80198 8296 80238 8336
rect 80238 8296 80263 8336
rect 80009 8273 80095 8296
rect 80177 8273 80263 8296
rect 95129 8336 95215 8359
rect 95297 8336 95383 8359
rect 95129 8296 95154 8336
rect 95154 8296 95194 8336
rect 95194 8296 95215 8336
rect 95297 8296 95318 8336
rect 95318 8296 95358 8336
rect 95358 8296 95383 8336
rect 95129 8273 95215 8296
rect 95297 8273 95383 8296
rect 3169 7580 3255 7603
rect 3337 7580 3423 7603
rect 3169 7540 3194 7580
rect 3194 7540 3234 7580
rect 3234 7540 3255 7580
rect 3337 7540 3358 7580
rect 3358 7540 3398 7580
rect 3398 7540 3423 7580
rect 3169 7517 3255 7540
rect 3337 7517 3423 7540
rect 18289 7580 18375 7603
rect 18457 7580 18543 7603
rect 18289 7540 18314 7580
rect 18314 7540 18354 7580
rect 18354 7540 18375 7580
rect 18457 7540 18478 7580
rect 18478 7540 18518 7580
rect 18518 7540 18543 7580
rect 18289 7517 18375 7540
rect 18457 7517 18543 7540
rect 33409 7580 33495 7603
rect 33577 7580 33663 7603
rect 33409 7540 33434 7580
rect 33434 7540 33474 7580
rect 33474 7540 33495 7580
rect 33577 7540 33598 7580
rect 33598 7540 33638 7580
rect 33638 7540 33663 7580
rect 33409 7517 33495 7540
rect 33577 7517 33663 7540
rect 48529 7580 48615 7603
rect 48697 7580 48783 7603
rect 48529 7540 48554 7580
rect 48554 7540 48594 7580
rect 48594 7540 48615 7580
rect 48697 7540 48718 7580
rect 48718 7540 48758 7580
rect 48758 7540 48783 7580
rect 48529 7517 48615 7540
rect 48697 7517 48783 7540
rect 63649 7580 63735 7603
rect 63817 7580 63903 7603
rect 63649 7540 63674 7580
rect 63674 7540 63714 7580
rect 63714 7540 63735 7580
rect 63817 7540 63838 7580
rect 63838 7540 63878 7580
rect 63878 7540 63903 7580
rect 63649 7517 63735 7540
rect 63817 7517 63903 7540
rect 78769 7580 78855 7603
rect 78937 7580 79023 7603
rect 78769 7540 78794 7580
rect 78794 7540 78834 7580
rect 78834 7540 78855 7580
rect 78937 7540 78958 7580
rect 78958 7540 78998 7580
rect 78998 7540 79023 7580
rect 78769 7517 78855 7540
rect 78937 7517 79023 7540
rect 93889 7580 93975 7603
rect 94057 7580 94143 7603
rect 93889 7540 93914 7580
rect 93914 7540 93954 7580
rect 93954 7540 93975 7580
rect 94057 7540 94078 7580
rect 94078 7540 94118 7580
rect 94118 7540 94143 7580
rect 93889 7517 93975 7540
rect 94057 7517 94143 7540
rect 4409 6824 4495 6847
rect 4577 6824 4663 6847
rect 4409 6784 4434 6824
rect 4434 6784 4474 6824
rect 4474 6784 4495 6824
rect 4577 6784 4598 6824
rect 4598 6784 4638 6824
rect 4638 6784 4663 6824
rect 4409 6761 4495 6784
rect 4577 6761 4663 6784
rect 19529 6824 19615 6847
rect 19697 6824 19783 6847
rect 19529 6784 19554 6824
rect 19554 6784 19594 6824
rect 19594 6784 19615 6824
rect 19697 6784 19718 6824
rect 19718 6784 19758 6824
rect 19758 6784 19783 6824
rect 19529 6761 19615 6784
rect 19697 6761 19783 6784
rect 34649 6824 34735 6847
rect 34817 6824 34903 6847
rect 34649 6784 34674 6824
rect 34674 6784 34714 6824
rect 34714 6784 34735 6824
rect 34817 6784 34838 6824
rect 34838 6784 34878 6824
rect 34878 6784 34903 6824
rect 34649 6761 34735 6784
rect 34817 6761 34903 6784
rect 49769 6824 49855 6847
rect 49937 6824 50023 6847
rect 49769 6784 49794 6824
rect 49794 6784 49834 6824
rect 49834 6784 49855 6824
rect 49937 6784 49958 6824
rect 49958 6784 49998 6824
rect 49998 6784 50023 6824
rect 49769 6761 49855 6784
rect 49937 6761 50023 6784
rect 64889 6824 64975 6847
rect 65057 6824 65143 6847
rect 64889 6784 64914 6824
rect 64914 6784 64954 6824
rect 64954 6784 64975 6824
rect 65057 6784 65078 6824
rect 65078 6784 65118 6824
rect 65118 6784 65143 6824
rect 64889 6761 64975 6784
rect 65057 6761 65143 6784
rect 80009 6824 80095 6847
rect 80177 6824 80263 6847
rect 80009 6784 80034 6824
rect 80034 6784 80074 6824
rect 80074 6784 80095 6824
rect 80177 6784 80198 6824
rect 80198 6784 80238 6824
rect 80238 6784 80263 6824
rect 80009 6761 80095 6784
rect 80177 6761 80263 6784
rect 95129 6824 95215 6847
rect 95297 6824 95383 6847
rect 95129 6784 95154 6824
rect 95154 6784 95194 6824
rect 95194 6784 95215 6824
rect 95297 6784 95318 6824
rect 95318 6784 95358 6824
rect 95358 6784 95383 6824
rect 95129 6761 95215 6784
rect 95297 6761 95383 6784
rect 3169 6068 3255 6091
rect 3337 6068 3423 6091
rect 3169 6028 3194 6068
rect 3194 6028 3234 6068
rect 3234 6028 3255 6068
rect 3337 6028 3358 6068
rect 3358 6028 3398 6068
rect 3398 6028 3423 6068
rect 3169 6005 3255 6028
rect 3337 6005 3423 6028
rect 18289 6068 18375 6091
rect 18457 6068 18543 6091
rect 18289 6028 18314 6068
rect 18314 6028 18354 6068
rect 18354 6028 18375 6068
rect 18457 6028 18478 6068
rect 18478 6028 18518 6068
rect 18518 6028 18543 6068
rect 18289 6005 18375 6028
rect 18457 6005 18543 6028
rect 33409 6068 33495 6091
rect 33577 6068 33663 6091
rect 33409 6028 33434 6068
rect 33434 6028 33474 6068
rect 33474 6028 33495 6068
rect 33577 6028 33598 6068
rect 33598 6028 33638 6068
rect 33638 6028 33663 6068
rect 33409 6005 33495 6028
rect 33577 6005 33663 6028
rect 48529 6068 48615 6091
rect 48697 6068 48783 6091
rect 48529 6028 48554 6068
rect 48554 6028 48594 6068
rect 48594 6028 48615 6068
rect 48697 6028 48718 6068
rect 48718 6028 48758 6068
rect 48758 6028 48783 6068
rect 48529 6005 48615 6028
rect 48697 6005 48783 6028
rect 63649 6068 63735 6091
rect 63817 6068 63903 6091
rect 63649 6028 63674 6068
rect 63674 6028 63714 6068
rect 63714 6028 63735 6068
rect 63817 6028 63838 6068
rect 63838 6028 63878 6068
rect 63878 6028 63903 6068
rect 63649 6005 63735 6028
rect 63817 6005 63903 6028
rect 78769 6068 78855 6091
rect 78937 6068 79023 6091
rect 78769 6028 78794 6068
rect 78794 6028 78834 6068
rect 78834 6028 78855 6068
rect 78937 6028 78958 6068
rect 78958 6028 78998 6068
rect 78998 6028 79023 6068
rect 78769 6005 78855 6028
rect 78937 6005 79023 6028
rect 93889 6068 93975 6091
rect 94057 6068 94143 6091
rect 93889 6028 93914 6068
rect 93914 6028 93954 6068
rect 93954 6028 93975 6068
rect 94057 6028 94078 6068
rect 94078 6028 94118 6068
rect 94118 6028 94143 6068
rect 93889 6005 93975 6028
rect 94057 6005 94143 6028
rect 4409 5312 4495 5335
rect 4577 5312 4663 5335
rect 4409 5272 4434 5312
rect 4434 5272 4474 5312
rect 4474 5272 4495 5312
rect 4577 5272 4598 5312
rect 4598 5272 4638 5312
rect 4638 5272 4663 5312
rect 4409 5249 4495 5272
rect 4577 5249 4663 5272
rect 19529 5312 19615 5335
rect 19697 5312 19783 5335
rect 19529 5272 19554 5312
rect 19554 5272 19594 5312
rect 19594 5272 19615 5312
rect 19697 5272 19718 5312
rect 19718 5272 19758 5312
rect 19758 5272 19783 5312
rect 19529 5249 19615 5272
rect 19697 5249 19783 5272
rect 34649 5312 34735 5335
rect 34817 5312 34903 5335
rect 34649 5272 34674 5312
rect 34674 5272 34714 5312
rect 34714 5272 34735 5312
rect 34817 5272 34838 5312
rect 34838 5272 34878 5312
rect 34878 5272 34903 5312
rect 34649 5249 34735 5272
rect 34817 5249 34903 5272
rect 49769 5312 49855 5335
rect 49937 5312 50023 5335
rect 49769 5272 49794 5312
rect 49794 5272 49834 5312
rect 49834 5272 49855 5312
rect 49937 5272 49958 5312
rect 49958 5272 49998 5312
rect 49998 5272 50023 5312
rect 49769 5249 49855 5272
rect 49937 5249 50023 5272
rect 64889 5312 64975 5335
rect 65057 5312 65143 5335
rect 64889 5272 64914 5312
rect 64914 5272 64954 5312
rect 64954 5272 64975 5312
rect 65057 5272 65078 5312
rect 65078 5272 65118 5312
rect 65118 5272 65143 5312
rect 64889 5249 64975 5272
rect 65057 5249 65143 5272
rect 80009 5312 80095 5335
rect 80177 5312 80263 5335
rect 80009 5272 80034 5312
rect 80034 5272 80074 5312
rect 80074 5272 80095 5312
rect 80177 5272 80198 5312
rect 80198 5272 80238 5312
rect 80238 5272 80263 5312
rect 80009 5249 80095 5272
rect 80177 5249 80263 5272
rect 95129 5312 95215 5335
rect 95297 5312 95383 5335
rect 95129 5272 95154 5312
rect 95154 5272 95194 5312
rect 95194 5272 95215 5312
rect 95297 5272 95318 5312
rect 95318 5272 95358 5312
rect 95358 5272 95383 5312
rect 95129 5249 95215 5272
rect 95297 5249 95383 5272
rect 3169 4556 3255 4579
rect 3337 4556 3423 4579
rect 3169 4516 3194 4556
rect 3194 4516 3234 4556
rect 3234 4516 3255 4556
rect 3337 4516 3358 4556
rect 3358 4516 3398 4556
rect 3398 4516 3423 4556
rect 3169 4493 3255 4516
rect 3337 4493 3423 4516
rect 18289 4556 18375 4579
rect 18457 4556 18543 4579
rect 18289 4516 18314 4556
rect 18314 4516 18354 4556
rect 18354 4516 18375 4556
rect 18457 4516 18478 4556
rect 18478 4516 18518 4556
rect 18518 4516 18543 4556
rect 18289 4493 18375 4516
rect 18457 4493 18543 4516
rect 33409 4556 33495 4579
rect 33577 4556 33663 4579
rect 33409 4516 33434 4556
rect 33434 4516 33474 4556
rect 33474 4516 33495 4556
rect 33577 4516 33598 4556
rect 33598 4516 33638 4556
rect 33638 4516 33663 4556
rect 33409 4493 33495 4516
rect 33577 4493 33663 4516
rect 48529 4556 48615 4579
rect 48697 4556 48783 4579
rect 48529 4516 48554 4556
rect 48554 4516 48594 4556
rect 48594 4516 48615 4556
rect 48697 4516 48718 4556
rect 48718 4516 48758 4556
rect 48758 4516 48783 4556
rect 48529 4493 48615 4516
rect 48697 4493 48783 4516
rect 63649 4556 63735 4579
rect 63817 4556 63903 4579
rect 63649 4516 63674 4556
rect 63674 4516 63714 4556
rect 63714 4516 63735 4556
rect 63817 4516 63838 4556
rect 63838 4516 63878 4556
rect 63878 4516 63903 4556
rect 63649 4493 63735 4516
rect 63817 4493 63903 4516
rect 78769 4556 78855 4579
rect 78937 4556 79023 4579
rect 78769 4516 78794 4556
rect 78794 4516 78834 4556
rect 78834 4516 78855 4556
rect 78937 4516 78958 4556
rect 78958 4516 78998 4556
rect 78998 4516 79023 4556
rect 78769 4493 78855 4516
rect 78937 4493 79023 4516
rect 93889 4556 93975 4579
rect 94057 4556 94143 4579
rect 93889 4516 93914 4556
rect 93914 4516 93954 4556
rect 93954 4516 93975 4556
rect 94057 4516 94078 4556
rect 94078 4516 94118 4556
rect 94118 4516 94143 4556
rect 93889 4493 93975 4516
rect 94057 4493 94143 4516
rect 4409 3800 4495 3823
rect 4577 3800 4663 3823
rect 4409 3760 4434 3800
rect 4434 3760 4474 3800
rect 4474 3760 4495 3800
rect 4577 3760 4598 3800
rect 4598 3760 4638 3800
rect 4638 3760 4663 3800
rect 4409 3737 4495 3760
rect 4577 3737 4663 3760
rect 19529 3800 19615 3823
rect 19697 3800 19783 3823
rect 19529 3760 19554 3800
rect 19554 3760 19594 3800
rect 19594 3760 19615 3800
rect 19697 3760 19718 3800
rect 19718 3760 19758 3800
rect 19758 3760 19783 3800
rect 19529 3737 19615 3760
rect 19697 3737 19783 3760
rect 34649 3800 34735 3823
rect 34817 3800 34903 3823
rect 34649 3760 34674 3800
rect 34674 3760 34714 3800
rect 34714 3760 34735 3800
rect 34817 3760 34838 3800
rect 34838 3760 34878 3800
rect 34878 3760 34903 3800
rect 34649 3737 34735 3760
rect 34817 3737 34903 3760
rect 49769 3800 49855 3823
rect 49937 3800 50023 3823
rect 49769 3760 49794 3800
rect 49794 3760 49834 3800
rect 49834 3760 49855 3800
rect 49937 3760 49958 3800
rect 49958 3760 49998 3800
rect 49998 3760 50023 3800
rect 49769 3737 49855 3760
rect 49937 3737 50023 3760
rect 64889 3800 64975 3823
rect 65057 3800 65143 3823
rect 64889 3760 64914 3800
rect 64914 3760 64954 3800
rect 64954 3760 64975 3800
rect 65057 3760 65078 3800
rect 65078 3760 65118 3800
rect 65118 3760 65143 3800
rect 64889 3737 64975 3760
rect 65057 3737 65143 3760
rect 80009 3800 80095 3823
rect 80177 3800 80263 3823
rect 80009 3760 80034 3800
rect 80034 3760 80074 3800
rect 80074 3760 80095 3800
rect 80177 3760 80198 3800
rect 80198 3760 80238 3800
rect 80238 3760 80263 3800
rect 80009 3737 80095 3760
rect 80177 3737 80263 3760
rect 95129 3800 95215 3823
rect 95297 3800 95383 3823
rect 95129 3760 95154 3800
rect 95154 3760 95194 3800
rect 95194 3760 95215 3800
rect 95297 3760 95318 3800
rect 95318 3760 95358 3800
rect 95358 3760 95383 3800
rect 95129 3737 95215 3760
rect 95297 3737 95383 3760
rect 3169 3044 3255 3067
rect 3337 3044 3423 3067
rect 3169 3004 3194 3044
rect 3194 3004 3234 3044
rect 3234 3004 3255 3044
rect 3337 3004 3358 3044
rect 3358 3004 3398 3044
rect 3398 3004 3423 3044
rect 3169 2981 3255 3004
rect 3337 2981 3423 3004
rect 18289 3044 18375 3067
rect 18457 3044 18543 3067
rect 18289 3004 18314 3044
rect 18314 3004 18354 3044
rect 18354 3004 18375 3044
rect 18457 3004 18478 3044
rect 18478 3004 18518 3044
rect 18518 3004 18543 3044
rect 18289 2981 18375 3004
rect 18457 2981 18543 3004
rect 33409 3044 33495 3067
rect 33577 3044 33663 3067
rect 33409 3004 33434 3044
rect 33434 3004 33474 3044
rect 33474 3004 33495 3044
rect 33577 3004 33598 3044
rect 33598 3004 33638 3044
rect 33638 3004 33663 3044
rect 33409 2981 33495 3004
rect 33577 2981 33663 3004
rect 48529 3044 48615 3067
rect 48697 3044 48783 3067
rect 48529 3004 48554 3044
rect 48554 3004 48594 3044
rect 48594 3004 48615 3044
rect 48697 3004 48718 3044
rect 48718 3004 48758 3044
rect 48758 3004 48783 3044
rect 48529 2981 48615 3004
rect 48697 2981 48783 3004
rect 63649 3044 63735 3067
rect 63817 3044 63903 3067
rect 63649 3004 63674 3044
rect 63674 3004 63714 3044
rect 63714 3004 63735 3044
rect 63817 3004 63838 3044
rect 63838 3004 63878 3044
rect 63878 3004 63903 3044
rect 63649 2981 63735 3004
rect 63817 2981 63903 3004
rect 78769 3044 78855 3067
rect 78937 3044 79023 3067
rect 78769 3004 78794 3044
rect 78794 3004 78834 3044
rect 78834 3004 78855 3044
rect 78937 3004 78958 3044
rect 78958 3004 78998 3044
rect 78998 3004 79023 3044
rect 78769 2981 78855 3004
rect 78937 2981 79023 3004
rect 93889 3044 93975 3067
rect 94057 3044 94143 3067
rect 93889 3004 93914 3044
rect 93914 3004 93954 3044
rect 93954 3004 93975 3044
rect 94057 3004 94078 3044
rect 94078 3004 94118 3044
rect 94118 3004 94143 3044
rect 93889 2981 93975 3004
rect 94057 2981 94143 3004
rect 4409 2288 4495 2311
rect 4577 2288 4663 2311
rect 4409 2248 4434 2288
rect 4434 2248 4474 2288
rect 4474 2248 4495 2288
rect 4577 2248 4598 2288
rect 4598 2248 4638 2288
rect 4638 2248 4663 2288
rect 4409 2225 4495 2248
rect 4577 2225 4663 2248
rect 19529 2288 19615 2311
rect 19697 2288 19783 2311
rect 19529 2248 19554 2288
rect 19554 2248 19594 2288
rect 19594 2248 19615 2288
rect 19697 2248 19718 2288
rect 19718 2248 19758 2288
rect 19758 2248 19783 2288
rect 19529 2225 19615 2248
rect 19697 2225 19783 2248
rect 34649 2288 34735 2311
rect 34817 2288 34903 2311
rect 34649 2248 34674 2288
rect 34674 2248 34714 2288
rect 34714 2248 34735 2288
rect 34817 2248 34838 2288
rect 34838 2248 34878 2288
rect 34878 2248 34903 2288
rect 34649 2225 34735 2248
rect 34817 2225 34903 2248
rect 49769 2288 49855 2311
rect 49937 2288 50023 2311
rect 49769 2248 49794 2288
rect 49794 2248 49834 2288
rect 49834 2248 49855 2288
rect 49937 2248 49958 2288
rect 49958 2248 49998 2288
rect 49998 2248 50023 2288
rect 49769 2225 49855 2248
rect 49937 2225 50023 2248
rect 64889 2288 64975 2311
rect 65057 2288 65143 2311
rect 64889 2248 64914 2288
rect 64914 2248 64954 2288
rect 64954 2248 64975 2288
rect 65057 2248 65078 2288
rect 65078 2248 65118 2288
rect 65118 2248 65143 2288
rect 64889 2225 64975 2248
rect 65057 2225 65143 2248
rect 80009 2288 80095 2311
rect 80177 2288 80263 2311
rect 80009 2248 80034 2288
rect 80034 2248 80074 2288
rect 80074 2248 80095 2288
rect 80177 2248 80198 2288
rect 80198 2248 80238 2288
rect 80238 2248 80263 2288
rect 80009 2225 80095 2248
rect 80177 2225 80263 2248
rect 95129 2288 95215 2311
rect 95297 2288 95383 2311
rect 95129 2248 95154 2288
rect 95154 2248 95194 2288
rect 95194 2248 95215 2288
rect 95297 2248 95318 2288
rect 95318 2248 95358 2288
rect 95358 2248 95383 2288
rect 95129 2225 95215 2248
rect 95297 2225 95383 2248
rect 3169 1532 3255 1555
rect 3337 1532 3423 1555
rect 3169 1492 3194 1532
rect 3194 1492 3234 1532
rect 3234 1492 3255 1532
rect 3337 1492 3358 1532
rect 3358 1492 3398 1532
rect 3398 1492 3423 1532
rect 3169 1469 3255 1492
rect 3337 1469 3423 1492
rect 18289 1532 18375 1555
rect 18457 1532 18543 1555
rect 18289 1492 18314 1532
rect 18314 1492 18354 1532
rect 18354 1492 18375 1532
rect 18457 1492 18478 1532
rect 18478 1492 18518 1532
rect 18518 1492 18543 1532
rect 18289 1469 18375 1492
rect 18457 1469 18543 1492
rect 33409 1532 33495 1555
rect 33577 1532 33663 1555
rect 33409 1492 33434 1532
rect 33434 1492 33474 1532
rect 33474 1492 33495 1532
rect 33577 1492 33598 1532
rect 33598 1492 33638 1532
rect 33638 1492 33663 1532
rect 33409 1469 33495 1492
rect 33577 1469 33663 1492
rect 48529 1532 48615 1555
rect 48697 1532 48783 1555
rect 48529 1492 48554 1532
rect 48554 1492 48594 1532
rect 48594 1492 48615 1532
rect 48697 1492 48718 1532
rect 48718 1492 48758 1532
rect 48758 1492 48783 1532
rect 48529 1469 48615 1492
rect 48697 1469 48783 1492
rect 63649 1532 63735 1555
rect 63817 1532 63903 1555
rect 63649 1492 63674 1532
rect 63674 1492 63714 1532
rect 63714 1492 63735 1532
rect 63817 1492 63838 1532
rect 63838 1492 63878 1532
rect 63878 1492 63903 1532
rect 63649 1469 63735 1492
rect 63817 1469 63903 1492
rect 78769 1532 78855 1555
rect 78937 1532 79023 1555
rect 78769 1492 78794 1532
rect 78794 1492 78834 1532
rect 78834 1492 78855 1532
rect 78937 1492 78958 1532
rect 78958 1492 78998 1532
rect 78998 1492 79023 1532
rect 78769 1469 78855 1492
rect 78937 1469 79023 1492
rect 93889 1532 93975 1555
rect 94057 1532 94143 1555
rect 93889 1492 93914 1532
rect 93914 1492 93954 1532
rect 93954 1492 93975 1532
rect 94057 1492 94078 1532
rect 94078 1492 94118 1532
rect 94118 1492 94143 1532
rect 93889 1469 93975 1492
rect 94057 1469 94143 1492
rect 4409 776 4495 799
rect 4577 776 4663 799
rect 4409 736 4434 776
rect 4434 736 4474 776
rect 4474 736 4495 776
rect 4577 736 4598 776
rect 4598 736 4638 776
rect 4638 736 4663 776
rect 4409 713 4495 736
rect 4577 713 4663 736
rect 19529 776 19615 799
rect 19697 776 19783 799
rect 19529 736 19554 776
rect 19554 736 19594 776
rect 19594 736 19615 776
rect 19697 736 19718 776
rect 19718 736 19758 776
rect 19758 736 19783 776
rect 19529 713 19615 736
rect 19697 713 19783 736
rect 34649 776 34735 799
rect 34817 776 34903 799
rect 34649 736 34674 776
rect 34674 736 34714 776
rect 34714 736 34735 776
rect 34817 736 34838 776
rect 34838 736 34878 776
rect 34878 736 34903 776
rect 34649 713 34735 736
rect 34817 713 34903 736
rect 49769 776 49855 799
rect 49937 776 50023 799
rect 49769 736 49794 776
rect 49794 736 49834 776
rect 49834 736 49855 776
rect 49937 736 49958 776
rect 49958 736 49998 776
rect 49998 736 50023 776
rect 49769 713 49855 736
rect 49937 713 50023 736
rect 64889 776 64975 799
rect 65057 776 65143 799
rect 64889 736 64914 776
rect 64914 736 64954 776
rect 64954 736 64975 776
rect 65057 736 65078 776
rect 65078 736 65118 776
rect 65118 736 65143 776
rect 64889 713 64975 736
rect 65057 713 65143 736
rect 80009 776 80095 799
rect 80177 776 80263 799
rect 80009 736 80034 776
rect 80034 736 80074 776
rect 80074 736 80095 776
rect 80177 736 80198 776
rect 80198 736 80238 776
rect 80238 736 80263 776
rect 80009 713 80095 736
rect 80177 713 80263 736
rect 95129 776 95215 799
rect 95297 776 95383 799
rect 95129 736 95154 776
rect 95154 736 95194 776
rect 95194 736 95215 776
rect 95297 736 95318 776
rect 95318 736 95358 776
rect 95358 736 95383 776
rect 95129 713 95215 736
rect 95297 713 95383 736
<< metal6 >>
rect 3076 37843 3516 38600
rect 3076 37757 3169 37843
rect 3255 37757 3337 37843
rect 3423 37757 3516 37843
rect 3076 36331 3516 37757
rect 3076 36245 3169 36331
rect 3255 36245 3337 36331
rect 3423 36245 3516 36331
rect 3076 34819 3516 36245
rect 3076 34733 3169 34819
rect 3255 34733 3337 34819
rect 3423 34733 3516 34819
rect 3076 33307 3516 34733
rect 3076 33221 3169 33307
rect 3255 33221 3337 33307
rect 3423 33221 3516 33307
rect 3076 31795 3516 33221
rect 3076 31709 3169 31795
rect 3255 31709 3337 31795
rect 3423 31709 3516 31795
rect 3076 30283 3516 31709
rect 3076 30197 3169 30283
rect 3255 30197 3337 30283
rect 3423 30197 3516 30283
rect 3076 28771 3516 30197
rect 3076 28685 3169 28771
rect 3255 28685 3337 28771
rect 3423 28685 3516 28771
rect 3076 27259 3516 28685
rect 3076 27173 3169 27259
rect 3255 27173 3337 27259
rect 3423 27173 3516 27259
rect 3076 25747 3516 27173
rect 3076 25661 3169 25747
rect 3255 25661 3337 25747
rect 3423 25661 3516 25747
rect 3076 24235 3516 25661
rect 3076 24149 3169 24235
rect 3255 24149 3337 24235
rect 3423 24149 3516 24235
rect 3076 22723 3516 24149
rect 3076 22637 3169 22723
rect 3255 22637 3337 22723
rect 3423 22637 3516 22723
rect 3076 21211 3516 22637
rect 3076 21125 3169 21211
rect 3255 21125 3337 21211
rect 3423 21125 3516 21211
rect 3076 19699 3516 21125
rect 3076 19613 3169 19699
rect 3255 19613 3337 19699
rect 3423 19613 3516 19699
rect 3076 18187 3516 19613
rect 3076 18101 3169 18187
rect 3255 18101 3337 18187
rect 3423 18101 3516 18187
rect 3076 16675 3516 18101
rect 3076 16589 3169 16675
rect 3255 16589 3337 16675
rect 3423 16589 3516 16675
rect 3076 15163 3516 16589
rect 3076 15077 3169 15163
rect 3255 15077 3337 15163
rect 3423 15077 3516 15163
rect 3076 13651 3516 15077
rect 3076 13565 3169 13651
rect 3255 13565 3337 13651
rect 3423 13565 3516 13651
rect 3076 12139 3516 13565
rect 3076 12053 3169 12139
rect 3255 12053 3337 12139
rect 3423 12053 3516 12139
rect 3076 10627 3516 12053
rect 3076 10541 3169 10627
rect 3255 10541 3337 10627
rect 3423 10541 3516 10627
rect 3076 9115 3516 10541
rect 3076 9029 3169 9115
rect 3255 9029 3337 9115
rect 3423 9029 3516 9115
rect 3076 7603 3516 9029
rect 3076 7517 3169 7603
rect 3255 7517 3337 7603
rect 3423 7517 3516 7603
rect 3076 6091 3516 7517
rect 3076 6005 3169 6091
rect 3255 6005 3337 6091
rect 3423 6005 3516 6091
rect 3076 4579 3516 6005
rect 3076 4493 3169 4579
rect 3255 4493 3337 4579
rect 3423 4493 3516 4579
rect 3076 3067 3516 4493
rect 3076 2981 3169 3067
rect 3255 2981 3337 3067
rect 3423 2981 3516 3067
rect 3076 1555 3516 2981
rect 3076 1469 3169 1555
rect 3255 1469 3337 1555
rect 3423 1469 3516 1555
rect 3076 712 3516 1469
rect 4316 38599 4756 38682
rect 4316 38513 4409 38599
rect 4495 38513 4577 38599
rect 4663 38513 4756 38599
rect 4316 37087 4756 38513
rect 4316 37001 4409 37087
rect 4495 37001 4577 37087
rect 4663 37001 4756 37087
rect 4316 35575 4756 37001
rect 4316 35489 4409 35575
rect 4495 35489 4577 35575
rect 4663 35489 4756 35575
rect 4316 34063 4756 35489
rect 4316 33977 4409 34063
rect 4495 33977 4577 34063
rect 4663 33977 4756 34063
rect 4316 32551 4756 33977
rect 4316 32465 4409 32551
rect 4495 32465 4577 32551
rect 4663 32465 4756 32551
rect 4316 31039 4756 32465
rect 4316 30953 4409 31039
rect 4495 30953 4577 31039
rect 4663 30953 4756 31039
rect 4316 29527 4756 30953
rect 4316 29441 4409 29527
rect 4495 29441 4577 29527
rect 4663 29441 4756 29527
rect 4316 28015 4756 29441
rect 4316 27929 4409 28015
rect 4495 27929 4577 28015
rect 4663 27929 4756 28015
rect 4316 26503 4756 27929
rect 4316 26417 4409 26503
rect 4495 26417 4577 26503
rect 4663 26417 4756 26503
rect 4316 24991 4756 26417
rect 4316 24905 4409 24991
rect 4495 24905 4577 24991
rect 4663 24905 4756 24991
rect 4316 23479 4756 24905
rect 4316 23393 4409 23479
rect 4495 23393 4577 23479
rect 4663 23393 4756 23479
rect 4316 21967 4756 23393
rect 4316 21881 4409 21967
rect 4495 21881 4577 21967
rect 4663 21881 4756 21967
rect 4316 20455 4756 21881
rect 4316 20369 4409 20455
rect 4495 20369 4577 20455
rect 4663 20369 4756 20455
rect 4316 18943 4756 20369
rect 4316 18857 4409 18943
rect 4495 18857 4577 18943
rect 4663 18857 4756 18943
rect 4316 17431 4756 18857
rect 4316 17345 4409 17431
rect 4495 17345 4577 17431
rect 4663 17345 4756 17431
rect 4316 15919 4756 17345
rect 4316 15833 4409 15919
rect 4495 15833 4577 15919
rect 4663 15833 4756 15919
rect 4316 14407 4756 15833
rect 4316 14321 4409 14407
rect 4495 14321 4577 14407
rect 4663 14321 4756 14407
rect 4316 12895 4756 14321
rect 4316 12809 4409 12895
rect 4495 12809 4577 12895
rect 4663 12809 4756 12895
rect 4316 11383 4756 12809
rect 4316 11297 4409 11383
rect 4495 11297 4577 11383
rect 4663 11297 4756 11383
rect 4316 9871 4756 11297
rect 4316 9785 4409 9871
rect 4495 9785 4577 9871
rect 4663 9785 4756 9871
rect 4316 8359 4756 9785
rect 4316 8273 4409 8359
rect 4495 8273 4577 8359
rect 4663 8273 4756 8359
rect 4316 6847 4756 8273
rect 4316 6761 4409 6847
rect 4495 6761 4577 6847
rect 4663 6761 4756 6847
rect 4316 5335 4756 6761
rect 4316 5249 4409 5335
rect 4495 5249 4577 5335
rect 4663 5249 4756 5335
rect 4316 3823 4756 5249
rect 4316 3737 4409 3823
rect 4495 3737 4577 3823
rect 4663 3737 4756 3823
rect 4316 2311 4756 3737
rect 4316 2225 4409 2311
rect 4495 2225 4577 2311
rect 4663 2225 4756 2311
rect 4316 799 4756 2225
rect 4316 713 4409 799
rect 4495 713 4577 799
rect 4663 713 4756 799
rect 4316 630 4756 713
rect 18196 37843 18636 38600
rect 18196 37757 18289 37843
rect 18375 37757 18457 37843
rect 18543 37757 18636 37843
rect 18196 36331 18636 37757
rect 18196 36245 18289 36331
rect 18375 36245 18457 36331
rect 18543 36245 18636 36331
rect 18196 34819 18636 36245
rect 18196 34733 18289 34819
rect 18375 34733 18457 34819
rect 18543 34733 18636 34819
rect 18196 33307 18636 34733
rect 18196 33221 18289 33307
rect 18375 33221 18457 33307
rect 18543 33221 18636 33307
rect 18196 31795 18636 33221
rect 18196 31709 18289 31795
rect 18375 31709 18457 31795
rect 18543 31709 18636 31795
rect 18196 30283 18636 31709
rect 18196 30197 18289 30283
rect 18375 30197 18457 30283
rect 18543 30197 18636 30283
rect 18196 28771 18636 30197
rect 18196 28685 18289 28771
rect 18375 28685 18457 28771
rect 18543 28685 18636 28771
rect 18196 27259 18636 28685
rect 18196 27173 18289 27259
rect 18375 27173 18457 27259
rect 18543 27173 18636 27259
rect 18196 25747 18636 27173
rect 18196 25661 18289 25747
rect 18375 25661 18457 25747
rect 18543 25661 18636 25747
rect 18196 24235 18636 25661
rect 18196 24149 18289 24235
rect 18375 24149 18457 24235
rect 18543 24149 18636 24235
rect 18196 22723 18636 24149
rect 18196 22637 18289 22723
rect 18375 22637 18457 22723
rect 18543 22637 18636 22723
rect 18196 21211 18636 22637
rect 18196 21125 18289 21211
rect 18375 21125 18457 21211
rect 18543 21125 18636 21211
rect 18196 19699 18636 21125
rect 18196 19613 18289 19699
rect 18375 19613 18457 19699
rect 18543 19613 18636 19699
rect 18196 18187 18636 19613
rect 18196 18101 18289 18187
rect 18375 18101 18457 18187
rect 18543 18101 18636 18187
rect 18196 16675 18636 18101
rect 18196 16589 18289 16675
rect 18375 16589 18457 16675
rect 18543 16589 18636 16675
rect 18196 15163 18636 16589
rect 18196 15077 18289 15163
rect 18375 15077 18457 15163
rect 18543 15077 18636 15163
rect 18196 13651 18636 15077
rect 18196 13565 18289 13651
rect 18375 13565 18457 13651
rect 18543 13565 18636 13651
rect 18196 12139 18636 13565
rect 18196 12053 18289 12139
rect 18375 12053 18457 12139
rect 18543 12053 18636 12139
rect 18196 10627 18636 12053
rect 18196 10541 18289 10627
rect 18375 10541 18457 10627
rect 18543 10541 18636 10627
rect 18196 9115 18636 10541
rect 18196 9029 18289 9115
rect 18375 9029 18457 9115
rect 18543 9029 18636 9115
rect 18196 7603 18636 9029
rect 18196 7517 18289 7603
rect 18375 7517 18457 7603
rect 18543 7517 18636 7603
rect 18196 6091 18636 7517
rect 18196 6005 18289 6091
rect 18375 6005 18457 6091
rect 18543 6005 18636 6091
rect 18196 4579 18636 6005
rect 18196 4493 18289 4579
rect 18375 4493 18457 4579
rect 18543 4493 18636 4579
rect 18196 3067 18636 4493
rect 18196 2981 18289 3067
rect 18375 2981 18457 3067
rect 18543 2981 18636 3067
rect 18196 1555 18636 2981
rect 18196 1469 18289 1555
rect 18375 1469 18457 1555
rect 18543 1469 18636 1555
rect 18196 712 18636 1469
rect 19436 38599 19876 38682
rect 19436 38513 19529 38599
rect 19615 38513 19697 38599
rect 19783 38513 19876 38599
rect 19436 37087 19876 38513
rect 19436 37001 19529 37087
rect 19615 37001 19697 37087
rect 19783 37001 19876 37087
rect 19436 35575 19876 37001
rect 19436 35489 19529 35575
rect 19615 35489 19697 35575
rect 19783 35489 19876 35575
rect 19436 34063 19876 35489
rect 19436 33977 19529 34063
rect 19615 33977 19697 34063
rect 19783 33977 19876 34063
rect 19436 32551 19876 33977
rect 19436 32465 19529 32551
rect 19615 32465 19697 32551
rect 19783 32465 19876 32551
rect 19436 31039 19876 32465
rect 19436 30953 19529 31039
rect 19615 30953 19697 31039
rect 19783 30953 19876 31039
rect 19436 29527 19876 30953
rect 19436 29441 19529 29527
rect 19615 29441 19697 29527
rect 19783 29441 19876 29527
rect 19436 28015 19876 29441
rect 19436 27929 19529 28015
rect 19615 27929 19697 28015
rect 19783 27929 19876 28015
rect 19436 26503 19876 27929
rect 19436 26417 19529 26503
rect 19615 26417 19697 26503
rect 19783 26417 19876 26503
rect 19436 24991 19876 26417
rect 19436 24905 19529 24991
rect 19615 24905 19697 24991
rect 19783 24905 19876 24991
rect 19436 23479 19876 24905
rect 19436 23393 19529 23479
rect 19615 23393 19697 23479
rect 19783 23393 19876 23479
rect 19436 21967 19876 23393
rect 19436 21881 19529 21967
rect 19615 21881 19697 21967
rect 19783 21881 19876 21967
rect 19436 20455 19876 21881
rect 19436 20369 19529 20455
rect 19615 20369 19697 20455
rect 19783 20369 19876 20455
rect 19436 18943 19876 20369
rect 19436 18857 19529 18943
rect 19615 18857 19697 18943
rect 19783 18857 19876 18943
rect 19436 17431 19876 18857
rect 19436 17345 19529 17431
rect 19615 17345 19697 17431
rect 19783 17345 19876 17431
rect 19436 15919 19876 17345
rect 19436 15833 19529 15919
rect 19615 15833 19697 15919
rect 19783 15833 19876 15919
rect 19436 14407 19876 15833
rect 19436 14321 19529 14407
rect 19615 14321 19697 14407
rect 19783 14321 19876 14407
rect 19436 12895 19876 14321
rect 19436 12809 19529 12895
rect 19615 12809 19697 12895
rect 19783 12809 19876 12895
rect 19436 11383 19876 12809
rect 19436 11297 19529 11383
rect 19615 11297 19697 11383
rect 19783 11297 19876 11383
rect 19436 9871 19876 11297
rect 19436 9785 19529 9871
rect 19615 9785 19697 9871
rect 19783 9785 19876 9871
rect 19436 8359 19876 9785
rect 19436 8273 19529 8359
rect 19615 8273 19697 8359
rect 19783 8273 19876 8359
rect 19436 6847 19876 8273
rect 19436 6761 19529 6847
rect 19615 6761 19697 6847
rect 19783 6761 19876 6847
rect 19436 5335 19876 6761
rect 19436 5249 19529 5335
rect 19615 5249 19697 5335
rect 19783 5249 19876 5335
rect 19436 3823 19876 5249
rect 19436 3737 19529 3823
rect 19615 3737 19697 3823
rect 19783 3737 19876 3823
rect 19436 2311 19876 3737
rect 19436 2225 19529 2311
rect 19615 2225 19697 2311
rect 19783 2225 19876 2311
rect 19436 799 19876 2225
rect 19436 713 19529 799
rect 19615 713 19697 799
rect 19783 713 19876 799
rect 19436 630 19876 713
rect 33316 37843 33756 38600
rect 33316 37757 33409 37843
rect 33495 37757 33577 37843
rect 33663 37757 33756 37843
rect 33316 36331 33756 37757
rect 33316 36245 33409 36331
rect 33495 36245 33577 36331
rect 33663 36245 33756 36331
rect 33316 34819 33756 36245
rect 33316 34733 33409 34819
rect 33495 34733 33577 34819
rect 33663 34733 33756 34819
rect 33316 33307 33756 34733
rect 33316 33221 33409 33307
rect 33495 33221 33577 33307
rect 33663 33221 33756 33307
rect 33316 31795 33756 33221
rect 33316 31709 33409 31795
rect 33495 31709 33577 31795
rect 33663 31709 33756 31795
rect 33316 30283 33756 31709
rect 33316 30197 33409 30283
rect 33495 30197 33577 30283
rect 33663 30197 33756 30283
rect 33316 28771 33756 30197
rect 33316 28685 33409 28771
rect 33495 28685 33577 28771
rect 33663 28685 33756 28771
rect 33316 27259 33756 28685
rect 33316 27173 33409 27259
rect 33495 27173 33577 27259
rect 33663 27173 33756 27259
rect 33316 25747 33756 27173
rect 33316 25661 33409 25747
rect 33495 25661 33577 25747
rect 33663 25661 33756 25747
rect 33316 24235 33756 25661
rect 33316 24149 33409 24235
rect 33495 24149 33577 24235
rect 33663 24149 33756 24235
rect 33316 22723 33756 24149
rect 33316 22637 33409 22723
rect 33495 22637 33577 22723
rect 33663 22637 33756 22723
rect 33316 21211 33756 22637
rect 33316 21125 33409 21211
rect 33495 21125 33577 21211
rect 33663 21125 33756 21211
rect 33316 19699 33756 21125
rect 33316 19613 33409 19699
rect 33495 19613 33577 19699
rect 33663 19613 33756 19699
rect 33316 18187 33756 19613
rect 33316 18101 33409 18187
rect 33495 18101 33577 18187
rect 33663 18101 33756 18187
rect 33316 16675 33756 18101
rect 33316 16589 33409 16675
rect 33495 16589 33577 16675
rect 33663 16589 33756 16675
rect 33316 15163 33756 16589
rect 33316 15077 33409 15163
rect 33495 15077 33577 15163
rect 33663 15077 33756 15163
rect 33316 13651 33756 15077
rect 33316 13565 33409 13651
rect 33495 13565 33577 13651
rect 33663 13565 33756 13651
rect 33316 12139 33756 13565
rect 33316 12053 33409 12139
rect 33495 12053 33577 12139
rect 33663 12053 33756 12139
rect 33316 10627 33756 12053
rect 33316 10541 33409 10627
rect 33495 10541 33577 10627
rect 33663 10541 33756 10627
rect 33316 9115 33756 10541
rect 33316 9029 33409 9115
rect 33495 9029 33577 9115
rect 33663 9029 33756 9115
rect 33316 7603 33756 9029
rect 33316 7517 33409 7603
rect 33495 7517 33577 7603
rect 33663 7517 33756 7603
rect 33316 6091 33756 7517
rect 33316 6005 33409 6091
rect 33495 6005 33577 6091
rect 33663 6005 33756 6091
rect 33316 4579 33756 6005
rect 33316 4493 33409 4579
rect 33495 4493 33577 4579
rect 33663 4493 33756 4579
rect 33316 3067 33756 4493
rect 33316 2981 33409 3067
rect 33495 2981 33577 3067
rect 33663 2981 33756 3067
rect 33316 1555 33756 2981
rect 33316 1469 33409 1555
rect 33495 1469 33577 1555
rect 33663 1469 33756 1555
rect 33316 712 33756 1469
rect 34556 38599 34996 38682
rect 34556 38513 34649 38599
rect 34735 38513 34817 38599
rect 34903 38513 34996 38599
rect 34556 37087 34996 38513
rect 34556 37001 34649 37087
rect 34735 37001 34817 37087
rect 34903 37001 34996 37087
rect 34556 35575 34996 37001
rect 34556 35489 34649 35575
rect 34735 35489 34817 35575
rect 34903 35489 34996 35575
rect 34556 34063 34996 35489
rect 34556 33977 34649 34063
rect 34735 33977 34817 34063
rect 34903 33977 34996 34063
rect 34556 32551 34996 33977
rect 34556 32465 34649 32551
rect 34735 32465 34817 32551
rect 34903 32465 34996 32551
rect 34556 31039 34996 32465
rect 34556 30953 34649 31039
rect 34735 30953 34817 31039
rect 34903 30953 34996 31039
rect 34556 29527 34996 30953
rect 34556 29441 34649 29527
rect 34735 29441 34817 29527
rect 34903 29441 34996 29527
rect 34556 28015 34996 29441
rect 34556 27929 34649 28015
rect 34735 27929 34817 28015
rect 34903 27929 34996 28015
rect 34556 26503 34996 27929
rect 34556 26417 34649 26503
rect 34735 26417 34817 26503
rect 34903 26417 34996 26503
rect 34556 24991 34996 26417
rect 34556 24905 34649 24991
rect 34735 24905 34817 24991
rect 34903 24905 34996 24991
rect 34556 23479 34996 24905
rect 34556 23393 34649 23479
rect 34735 23393 34817 23479
rect 34903 23393 34996 23479
rect 34556 21967 34996 23393
rect 34556 21881 34649 21967
rect 34735 21881 34817 21967
rect 34903 21881 34996 21967
rect 34556 20455 34996 21881
rect 34556 20369 34649 20455
rect 34735 20369 34817 20455
rect 34903 20369 34996 20455
rect 34556 18943 34996 20369
rect 34556 18857 34649 18943
rect 34735 18857 34817 18943
rect 34903 18857 34996 18943
rect 34556 17431 34996 18857
rect 34556 17345 34649 17431
rect 34735 17345 34817 17431
rect 34903 17345 34996 17431
rect 34556 15919 34996 17345
rect 34556 15833 34649 15919
rect 34735 15833 34817 15919
rect 34903 15833 34996 15919
rect 34556 14407 34996 15833
rect 34556 14321 34649 14407
rect 34735 14321 34817 14407
rect 34903 14321 34996 14407
rect 34556 12895 34996 14321
rect 34556 12809 34649 12895
rect 34735 12809 34817 12895
rect 34903 12809 34996 12895
rect 34556 11383 34996 12809
rect 34556 11297 34649 11383
rect 34735 11297 34817 11383
rect 34903 11297 34996 11383
rect 34556 9871 34996 11297
rect 34556 9785 34649 9871
rect 34735 9785 34817 9871
rect 34903 9785 34996 9871
rect 34556 8359 34996 9785
rect 34556 8273 34649 8359
rect 34735 8273 34817 8359
rect 34903 8273 34996 8359
rect 34556 6847 34996 8273
rect 34556 6761 34649 6847
rect 34735 6761 34817 6847
rect 34903 6761 34996 6847
rect 34556 5335 34996 6761
rect 34556 5249 34649 5335
rect 34735 5249 34817 5335
rect 34903 5249 34996 5335
rect 34556 3823 34996 5249
rect 34556 3737 34649 3823
rect 34735 3737 34817 3823
rect 34903 3737 34996 3823
rect 34556 2311 34996 3737
rect 34556 2225 34649 2311
rect 34735 2225 34817 2311
rect 34903 2225 34996 2311
rect 34556 799 34996 2225
rect 34556 713 34649 799
rect 34735 713 34817 799
rect 34903 713 34996 799
rect 34556 630 34996 713
rect 48436 37843 48876 38600
rect 48436 37757 48529 37843
rect 48615 37757 48697 37843
rect 48783 37757 48876 37843
rect 48436 36331 48876 37757
rect 48436 36245 48529 36331
rect 48615 36245 48697 36331
rect 48783 36245 48876 36331
rect 48436 34819 48876 36245
rect 48436 34733 48529 34819
rect 48615 34733 48697 34819
rect 48783 34733 48876 34819
rect 48436 33307 48876 34733
rect 48436 33221 48529 33307
rect 48615 33221 48697 33307
rect 48783 33221 48876 33307
rect 48436 31795 48876 33221
rect 48436 31709 48529 31795
rect 48615 31709 48697 31795
rect 48783 31709 48876 31795
rect 48436 30283 48876 31709
rect 48436 30197 48529 30283
rect 48615 30197 48697 30283
rect 48783 30197 48876 30283
rect 48436 28771 48876 30197
rect 48436 28685 48529 28771
rect 48615 28685 48697 28771
rect 48783 28685 48876 28771
rect 48436 27259 48876 28685
rect 48436 27173 48529 27259
rect 48615 27173 48697 27259
rect 48783 27173 48876 27259
rect 48436 25747 48876 27173
rect 48436 25661 48529 25747
rect 48615 25661 48697 25747
rect 48783 25661 48876 25747
rect 48436 24235 48876 25661
rect 48436 24149 48529 24235
rect 48615 24149 48697 24235
rect 48783 24149 48876 24235
rect 48436 22723 48876 24149
rect 48436 22637 48529 22723
rect 48615 22637 48697 22723
rect 48783 22637 48876 22723
rect 48436 21211 48876 22637
rect 48436 21125 48529 21211
rect 48615 21125 48697 21211
rect 48783 21125 48876 21211
rect 48436 19699 48876 21125
rect 48436 19613 48529 19699
rect 48615 19613 48697 19699
rect 48783 19613 48876 19699
rect 48436 18187 48876 19613
rect 48436 18101 48529 18187
rect 48615 18101 48697 18187
rect 48783 18101 48876 18187
rect 48436 16675 48876 18101
rect 48436 16589 48529 16675
rect 48615 16589 48697 16675
rect 48783 16589 48876 16675
rect 48436 15163 48876 16589
rect 48436 15077 48529 15163
rect 48615 15077 48697 15163
rect 48783 15077 48876 15163
rect 48436 13651 48876 15077
rect 48436 13565 48529 13651
rect 48615 13565 48697 13651
rect 48783 13565 48876 13651
rect 48436 12139 48876 13565
rect 48436 12053 48529 12139
rect 48615 12053 48697 12139
rect 48783 12053 48876 12139
rect 48436 10627 48876 12053
rect 48436 10541 48529 10627
rect 48615 10541 48697 10627
rect 48783 10541 48876 10627
rect 48436 9115 48876 10541
rect 48436 9029 48529 9115
rect 48615 9029 48697 9115
rect 48783 9029 48876 9115
rect 48436 7603 48876 9029
rect 48436 7517 48529 7603
rect 48615 7517 48697 7603
rect 48783 7517 48876 7603
rect 48436 6091 48876 7517
rect 48436 6005 48529 6091
rect 48615 6005 48697 6091
rect 48783 6005 48876 6091
rect 48436 4579 48876 6005
rect 48436 4493 48529 4579
rect 48615 4493 48697 4579
rect 48783 4493 48876 4579
rect 48436 3067 48876 4493
rect 48436 2981 48529 3067
rect 48615 2981 48697 3067
rect 48783 2981 48876 3067
rect 48436 1555 48876 2981
rect 48436 1469 48529 1555
rect 48615 1469 48697 1555
rect 48783 1469 48876 1555
rect 48436 712 48876 1469
rect 49676 38599 50116 38682
rect 49676 38513 49769 38599
rect 49855 38513 49937 38599
rect 50023 38513 50116 38599
rect 49676 37087 50116 38513
rect 49676 37001 49769 37087
rect 49855 37001 49937 37087
rect 50023 37001 50116 37087
rect 49676 35575 50116 37001
rect 49676 35489 49769 35575
rect 49855 35489 49937 35575
rect 50023 35489 50116 35575
rect 49676 34063 50116 35489
rect 49676 33977 49769 34063
rect 49855 33977 49937 34063
rect 50023 33977 50116 34063
rect 49676 32551 50116 33977
rect 49676 32465 49769 32551
rect 49855 32465 49937 32551
rect 50023 32465 50116 32551
rect 49676 31039 50116 32465
rect 49676 30953 49769 31039
rect 49855 30953 49937 31039
rect 50023 30953 50116 31039
rect 49676 29527 50116 30953
rect 49676 29441 49769 29527
rect 49855 29441 49937 29527
rect 50023 29441 50116 29527
rect 49676 28015 50116 29441
rect 49676 27929 49769 28015
rect 49855 27929 49937 28015
rect 50023 27929 50116 28015
rect 49676 26503 50116 27929
rect 49676 26417 49769 26503
rect 49855 26417 49937 26503
rect 50023 26417 50116 26503
rect 49676 24991 50116 26417
rect 49676 24905 49769 24991
rect 49855 24905 49937 24991
rect 50023 24905 50116 24991
rect 49676 23479 50116 24905
rect 49676 23393 49769 23479
rect 49855 23393 49937 23479
rect 50023 23393 50116 23479
rect 49676 21967 50116 23393
rect 49676 21881 49769 21967
rect 49855 21881 49937 21967
rect 50023 21881 50116 21967
rect 49676 20455 50116 21881
rect 49676 20369 49769 20455
rect 49855 20369 49937 20455
rect 50023 20369 50116 20455
rect 49676 18943 50116 20369
rect 49676 18857 49769 18943
rect 49855 18857 49937 18943
rect 50023 18857 50116 18943
rect 49676 17431 50116 18857
rect 49676 17345 49769 17431
rect 49855 17345 49937 17431
rect 50023 17345 50116 17431
rect 49676 15919 50116 17345
rect 49676 15833 49769 15919
rect 49855 15833 49937 15919
rect 50023 15833 50116 15919
rect 49676 14407 50116 15833
rect 49676 14321 49769 14407
rect 49855 14321 49937 14407
rect 50023 14321 50116 14407
rect 49676 12895 50116 14321
rect 49676 12809 49769 12895
rect 49855 12809 49937 12895
rect 50023 12809 50116 12895
rect 49676 11383 50116 12809
rect 49676 11297 49769 11383
rect 49855 11297 49937 11383
rect 50023 11297 50116 11383
rect 49676 9871 50116 11297
rect 49676 9785 49769 9871
rect 49855 9785 49937 9871
rect 50023 9785 50116 9871
rect 49676 8359 50116 9785
rect 49676 8273 49769 8359
rect 49855 8273 49937 8359
rect 50023 8273 50116 8359
rect 49676 6847 50116 8273
rect 49676 6761 49769 6847
rect 49855 6761 49937 6847
rect 50023 6761 50116 6847
rect 49676 5335 50116 6761
rect 49676 5249 49769 5335
rect 49855 5249 49937 5335
rect 50023 5249 50116 5335
rect 49676 3823 50116 5249
rect 49676 3737 49769 3823
rect 49855 3737 49937 3823
rect 50023 3737 50116 3823
rect 49676 2311 50116 3737
rect 49676 2225 49769 2311
rect 49855 2225 49937 2311
rect 50023 2225 50116 2311
rect 49676 799 50116 2225
rect 49676 713 49769 799
rect 49855 713 49937 799
rect 50023 713 50116 799
rect 49676 630 50116 713
rect 63556 37843 63996 38600
rect 63556 37757 63649 37843
rect 63735 37757 63817 37843
rect 63903 37757 63996 37843
rect 63556 36331 63996 37757
rect 63556 36245 63649 36331
rect 63735 36245 63817 36331
rect 63903 36245 63996 36331
rect 63556 34819 63996 36245
rect 63556 34733 63649 34819
rect 63735 34733 63817 34819
rect 63903 34733 63996 34819
rect 63556 33307 63996 34733
rect 63556 33221 63649 33307
rect 63735 33221 63817 33307
rect 63903 33221 63996 33307
rect 63556 31795 63996 33221
rect 63556 31709 63649 31795
rect 63735 31709 63817 31795
rect 63903 31709 63996 31795
rect 63556 30283 63996 31709
rect 63556 30197 63649 30283
rect 63735 30197 63817 30283
rect 63903 30197 63996 30283
rect 63556 28771 63996 30197
rect 63556 28685 63649 28771
rect 63735 28685 63817 28771
rect 63903 28685 63996 28771
rect 63556 27259 63996 28685
rect 63556 27173 63649 27259
rect 63735 27173 63817 27259
rect 63903 27173 63996 27259
rect 63556 25747 63996 27173
rect 63556 25661 63649 25747
rect 63735 25661 63817 25747
rect 63903 25661 63996 25747
rect 63556 24235 63996 25661
rect 63556 24149 63649 24235
rect 63735 24149 63817 24235
rect 63903 24149 63996 24235
rect 63556 22723 63996 24149
rect 63556 22637 63649 22723
rect 63735 22637 63817 22723
rect 63903 22637 63996 22723
rect 63556 21211 63996 22637
rect 63556 21125 63649 21211
rect 63735 21125 63817 21211
rect 63903 21125 63996 21211
rect 63556 19699 63996 21125
rect 63556 19613 63649 19699
rect 63735 19613 63817 19699
rect 63903 19613 63996 19699
rect 63556 18187 63996 19613
rect 63556 18101 63649 18187
rect 63735 18101 63817 18187
rect 63903 18101 63996 18187
rect 63556 16675 63996 18101
rect 63556 16589 63649 16675
rect 63735 16589 63817 16675
rect 63903 16589 63996 16675
rect 63556 15163 63996 16589
rect 63556 15077 63649 15163
rect 63735 15077 63817 15163
rect 63903 15077 63996 15163
rect 63556 13651 63996 15077
rect 63556 13565 63649 13651
rect 63735 13565 63817 13651
rect 63903 13565 63996 13651
rect 63556 12139 63996 13565
rect 63556 12053 63649 12139
rect 63735 12053 63817 12139
rect 63903 12053 63996 12139
rect 63556 10627 63996 12053
rect 63556 10541 63649 10627
rect 63735 10541 63817 10627
rect 63903 10541 63996 10627
rect 63556 9115 63996 10541
rect 63556 9029 63649 9115
rect 63735 9029 63817 9115
rect 63903 9029 63996 9115
rect 63556 7603 63996 9029
rect 63556 7517 63649 7603
rect 63735 7517 63817 7603
rect 63903 7517 63996 7603
rect 63556 6091 63996 7517
rect 63556 6005 63649 6091
rect 63735 6005 63817 6091
rect 63903 6005 63996 6091
rect 63556 4579 63996 6005
rect 63556 4493 63649 4579
rect 63735 4493 63817 4579
rect 63903 4493 63996 4579
rect 63556 3067 63996 4493
rect 63556 2981 63649 3067
rect 63735 2981 63817 3067
rect 63903 2981 63996 3067
rect 63556 1555 63996 2981
rect 63556 1469 63649 1555
rect 63735 1469 63817 1555
rect 63903 1469 63996 1555
rect 63556 712 63996 1469
rect 64796 38599 65236 38682
rect 64796 38513 64889 38599
rect 64975 38513 65057 38599
rect 65143 38513 65236 38599
rect 64796 37087 65236 38513
rect 64796 37001 64889 37087
rect 64975 37001 65057 37087
rect 65143 37001 65236 37087
rect 64796 35575 65236 37001
rect 64796 35489 64889 35575
rect 64975 35489 65057 35575
rect 65143 35489 65236 35575
rect 64796 34063 65236 35489
rect 64796 33977 64889 34063
rect 64975 33977 65057 34063
rect 65143 33977 65236 34063
rect 64796 32551 65236 33977
rect 64796 32465 64889 32551
rect 64975 32465 65057 32551
rect 65143 32465 65236 32551
rect 64796 31039 65236 32465
rect 64796 30953 64889 31039
rect 64975 30953 65057 31039
rect 65143 30953 65236 31039
rect 64796 29527 65236 30953
rect 64796 29441 64889 29527
rect 64975 29441 65057 29527
rect 65143 29441 65236 29527
rect 64796 28015 65236 29441
rect 64796 27929 64889 28015
rect 64975 27929 65057 28015
rect 65143 27929 65236 28015
rect 64796 26503 65236 27929
rect 64796 26417 64889 26503
rect 64975 26417 65057 26503
rect 65143 26417 65236 26503
rect 64796 24991 65236 26417
rect 64796 24905 64889 24991
rect 64975 24905 65057 24991
rect 65143 24905 65236 24991
rect 64796 23479 65236 24905
rect 64796 23393 64889 23479
rect 64975 23393 65057 23479
rect 65143 23393 65236 23479
rect 64796 21967 65236 23393
rect 64796 21881 64889 21967
rect 64975 21881 65057 21967
rect 65143 21881 65236 21967
rect 64796 20455 65236 21881
rect 64796 20369 64889 20455
rect 64975 20369 65057 20455
rect 65143 20369 65236 20455
rect 64796 18943 65236 20369
rect 64796 18857 64889 18943
rect 64975 18857 65057 18943
rect 65143 18857 65236 18943
rect 64796 17431 65236 18857
rect 64796 17345 64889 17431
rect 64975 17345 65057 17431
rect 65143 17345 65236 17431
rect 64796 15919 65236 17345
rect 64796 15833 64889 15919
rect 64975 15833 65057 15919
rect 65143 15833 65236 15919
rect 64796 14407 65236 15833
rect 64796 14321 64889 14407
rect 64975 14321 65057 14407
rect 65143 14321 65236 14407
rect 64796 12895 65236 14321
rect 64796 12809 64889 12895
rect 64975 12809 65057 12895
rect 65143 12809 65236 12895
rect 64796 11383 65236 12809
rect 64796 11297 64889 11383
rect 64975 11297 65057 11383
rect 65143 11297 65236 11383
rect 64796 9871 65236 11297
rect 64796 9785 64889 9871
rect 64975 9785 65057 9871
rect 65143 9785 65236 9871
rect 64796 8359 65236 9785
rect 64796 8273 64889 8359
rect 64975 8273 65057 8359
rect 65143 8273 65236 8359
rect 64796 6847 65236 8273
rect 64796 6761 64889 6847
rect 64975 6761 65057 6847
rect 65143 6761 65236 6847
rect 64796 5335 65236 6761
rect 64796 5249 64889 5335
rect 64975 5249 65057 5335
rect 65143 5249 65236 5335
rect 64796 3823 65236 5249
rect 64796 3737 64889 3823
rect 64975 3737 65057 3823
rect 65143 3737 65236 3823
rect 64796 2311 65236 3737
rect 64796 2225 64889 2311
rect 64975 2225 65057 2311
rect 65143 2225 65236 2311
rect 64796 799 65236 2225
rect 64796 713 64889 799
rect 64975 713 65057 799
rect 65143 713 65236 799
rect 64796 630 65236 713
rect 78676 37843 79116 38600
rect 78676 37757 78769 37843
rect 78855 37757 78937 37843
rect 79023 37757 79116 37843
rect 78676 36331 79116 37757
rect 78676 36245 78769 36331
rect 78855 36245 78937 36331
rect 79023 36245 79116 36331
rect 78676 34819 79116 36245
rect 78676 34733 78769 34819
rect 78855 34733 78937 34819
rect 79023 34733 79116 34819
rect 78676 33307 79116 34733
rect 78676 33221 78769 33307
rect 78855 33221 78937 33307
rect 79023 33221 79116 33307
rect 78676 31795 79116 33221
rect 78676 31709 78769 31795
rect 78855 31709 78937 31795
rect 79023 31709 79116 31795
rect 78676 30283 79116 31709
rect 78676 30197 78769 30283
rect 78855 30197 78937 30283
rect 79023 30197 79116 30283
rect 78676 28771 79116 30197
rect 78676 28685 78769 28771
rect 78855 28685 78937 28771
rect 79023 28685 79116 28771
rect 78676 27259 79116 28685
rect 78676 27173 78769 27259
rect 78855 27173 78937 27259
rect 79023 27173 79116 27259
rect 78676 25747 79116 27173
rect 78676 25661 78769 25747
rect 78855 25661 78937 25747
rect 79023 25661 79116 25747
rect 78676 24235 79116 25661
rect 78676 24149 78769 24235
rect 78855 24149 78937 24235
rect 79023 24149 79116 24235
rect 78676 22723 79116 24149
rect 78676 22637 78769 22723
rect 78855 22637 78937 22723
rect 79023 22637 79116 22723
rect 78676 21211 79116 22637
rect 78676 21125 78769 21211
rect 78855 21125 78937 21211
rect 79023 21125 79116 21211
rect 78676 19699 79116 21125
rect 78676 19613 78769 19699
rect 78855 19613 78937 19699
rect 79023 19613 79116 19699
rect 78676 18187 79116 19613
rect 78676 18101 78769 18187
rect 78855 18101 78937 18187
rect 79023 18101 79116 18187
rect 78676 16675 79116 18101
rect 78676 16589 78769 16675
rect 78855 16589 78937 16675
rect 79023 16589 79116 16675
rect 78676 15163 79116 16589
rect 78676 15077 78769 15163
rect 78855 15077 78937 15163
rect 79023 15077 79116 15163
rect 78676 13651 79116 15077
rect 78676 13565 78769 13651
rect 78855 13565 78937 13651
rect 79023 13565 79116 13651
rect 78676 12139 79116 13565
rect 78676 12053 78769 12139
rect 78855 12053 78937 12139
rect 79023 12053 79116 12139
rect 78676 10627 79116 12053
rect 78676 10541 78769 10627
rect 78855 10541 78937 10627
rect 79023 10541 79116 10627
rect 78676 9115 79116 10541
rect 78676 9029 78769 9115
rect 78855 9029 78937 9115
rect 79023 9029 79116 9115
rect 78676 7603 79116 9029
rect 78676 7517 78769 7603
rect 78855 7517 78937 7603
rect 79023 7517 79116 7603
rect 78676 6091 79116 7517
rect 78676 6005 78769 6091
rect 78855 6005 78937 6091
rect 79023 6005 79116 6091
rect 78676 4579 79116 6005
rect 78676 4493 78769 4579
rect 78855 4493 78937 4579
rect 79023 4493 79116 4579
rect 78676 3067 79116 4493
rect 78676 2981 78769 3067
rect 78855 2981 78937 3067
rect 79023 2981 79116 3067
rect 78676 1555 79116 2981
rect 78676 1469 78769 1555
rect 78855 1469 78937 1555
rect 79023 1469 79116 1555
rect 78676 712 79116 1469
rect 79916 38599 80356 38682
rect 79916 38513 80009 38599
rect 80095 38513 80177 38599
rect 80263 38513 80356 38599
rect 79916 37087 80356 38513
rect 79916 37001 80009 37087
rect 80095 37001 80177 37087
rect 80263 37001 80356 37087
rect 79916 35575 80356 37001
rect 79916 35489 80009 35575
rect 80095 35489 80177 35575
rect 80263 35489 80356 35575
rect 79916 34063 80356 35489
rect 79916 33977 80009 34063
rect 80095 33977 80177 34063
rect 80263 33977 80356 34063
rect 79916 32551 80356 33977
rect 79916 32465 80009 32551
rect 80095 32465 80177 32551
rect 80263 32465 80356 32551
rect 79916 31039 80356 32465
rect 79916 30953 80009 31039
rect 80095 30953 80177 31039
rect 80263 30953 80356 31039
rect 79916 29527 80356 30953
rect 79916 29441 80009 29527
rect 80095 29441 80177 29527
rect 80263 29441 80356 29527
rect 79916 28015 80356 29441
rect 79916 27929 80009 28015
rect 80095 27929 80177 28015
rect 80263 27929 80356 28015
rect 79916 26503 80356 27929
rect 79916 26417 80009 26503
rect 80095 26417 80177 26503
rect 80263 26417 80356 26503
rect 79916 24991 80356 26417
rect 79916 24905 80009 24991
rect 80095 24905 80177 24991
rect 80263 24905 80356 24991
rect 79916 23479 80356 24905
rect 79916 23393 80009 23479
rect 80095 23393 80177 23479
rect 80263 23393 80356 23479
rect 79916 21967 80356 23393
rect 79916 21881 80009 21967
rect 80095 21881 80177 21967
rect 80263 21881 80356 21967
rect 79916 20455 80356 21881
rect 79916 20369 80009 20455
rect 80095 20369 80177 20455
rect 80263 20369 80356 20455
rect 79916 18943 80356 20369
rect 79916 18857 80009 18943
rect 80095 18857 80177 18943
rect 80263 18857 80356 18943
rect 79916 17431 80356 18857
rect 79916 17345 80009 17431
rect 80095 17345 80177 17431
rect 80263 17345 80356 17431
rect 79916 15919 80356 17345
rect 79916 15833 80009 15919
rect 80095 15833 80177 15919
rect 80263 15833 80356 15919
rect 79916 14407 80356 15833
rect 79916 14321 80009 14407
rect 80095 14321 80177 14407
rect 80263 14321 80356 14407
rect 79916 12895 80356 14321
rect 79916 12809 80009 12895
rect 80095 12809 80177 12895
rect 80263 12809 80356 12895
rect 79916 11383 80356 12809
rect 79916 11297 80009 11383
rect 80095 11297 80177 11383
rect 80263 11297 80356 11383
rect 79916 9871 80356 11297
rect 79916 9785 80009 9871
rect 80095 9785 80177 9871
rect 80263 9785 80356 9871
rect 79916 8359 80356 9785
rect 79916 8273 80009 8359
rect 80095 8273 80177 8359
rect 80263 8273 80356 8359
rect 79916 6847 80356 8273
rect 79916 6761 80009 6847
rect 80095 6761 80177 6847
rect 80263 6761 80356 6847
rect 79916 5335 80356 6761
rect 79916 5249 80009 5335
rect 80095 5249 80177 5335
rect 80263 5249 80356 5335
rect 79916 3823 80356 5249
rect 79916 3737 80009 3823
rect 80095 3737 80177 3823
rect 80263 3737 80356 3823
rect 79916 2311 80356 3737
rect 79916 2225 80009 2311
rect 80095 2225 80177 2311
rect 80263 2225 80356 2311
rect 79916 799 80356 2225
rect 79916 713 80009 799
rect 80095 713 80177 799
rect 80263 713 80356 799
rect 79916 630 80356 713
rect 93796 37843 94236 38600
rect 93796 37757 93889 37843
rect 93975 37757 94057 37843
rect 94143 37757 94236 37843
rect 93796 36331 94236 37757
rect 93796 36245 93889 36331
rect 93975 36245 94057 36331
rect 94143 36245 94236 36331
rect 93796 34819 94236 36245
rect 93796 34733 93889 34819
rect 93975 34733 94057 34819
rect 94143 34733 94236 34819
rect 93796 33307 94236 34733
rect 93796 33221 93889 33307
rect 93975 33221 94057 33307
rect 94143 33221 94236 33307
rect 93796 31795 94236 33221
rect 93796 31709 93889 31795
rect 93975 31709 94057 31795
rect 94143 31709 94236 31795
rect 93796 30283 94236 31709
rect 93796 30197 93889 30283
rect 93975 30197 94057 30283
rect 94143 30197 94236 30283
rect 93796 28771 94236 30197
rect 93796 28685 93889 28771
rect 93975 28685 94057 28771
rect 94143 28685 94236 28771
rect 93796 27259 94236 28685
rect 93796 27173 93889 27259
rect 93975 27173 94057 27259
rect 94143 27173 94236 27259
rect 93796 25747 94236 27173
rect 93796 25661 93889 25747
rect 93975 25661 94057 25747
rect 94143 25661 94236 25747
rect 93796 24235 94236 25661
rect 93796 24149 93889 24235
rect 93975 24149 94057 24235
rect 94143 24149 94236 24235
rect 93796 22723 94236 24149
rect 93796 22637 93889 22723
rect 93975 22637 94057 22723
rect 94143 22637 94236 22723
rect 93796 21211 94236 22637
rect 93796 21125 93889 21211
rect 93975 21125 94057 21211
rect 94143 21125 94236 21211
rect 93796 19699 94236 21125
rect 93796 19613 93889 19699
rect 93975 19613 94057 19699
rect 94143 19613 94236 19699
rect 93796 18187 94236 19613
rect 93796 18101 93889 18187
rect 93975 18101 94057 18187
rect 94143 18101 94236 18187
rect 93796 16675 94236 18101
rect 93796 16589 93889 16675
rect 93975 16589 94057 16675
rect 94143 16589 94236 16675
rect 93796 15163 94236 16589
rect 93796 15077 93889 15163
rect 93975 15077 94057 15163
rect 94143 15077 94236 15163
rect 93796 13651 94236 15077
rect 93796 13565 93889 13651
rect 93975 13565 94057 13651
rect 94143 13565 94236 13651
rect 93796 12139 94236 13565
rect 93796 12053 93889 12139
rect 93975 12053 94057 12139
rect 94143 12053 94236 12139
rect 93796 10627 94236 12053
rect 93796 10541 93889 10627
rect 93975 10541 94057 10627
rect 94143 10541 94236 10627
rect 93796 9115 94236 10541
rect 93796 9029 93889 9115
rect 93975 9029 94057 9115
rect 94143 9029 94236 9115
rect 93796 7603 94236 9029
rect 93796 7517 93889 7603
rect 93975 7517 94057 7603
rect 94143 7517 94236 7603
rect 93796 6091 94236 7517
rect 93796 6005 93889 6091
rect 93975 6005 94057 6091
rect 94143 6005 94236 6091
rect 93796 4579 94236 6005
rect 93796 4493 93889 4579
rect 93975 4493 94057 4579
rect 94143 4493 94236 4579
rect 93796 3067 94236 4493
rect 93796 2981 93889 3067
rect 93975 2981 94057 3067
rect 94143 2981 94236 3067
rect 93796 1555 94236 2981
rect 93796 1469 93889 1555
rect 93975 1469 94057 1555
rect 94143 1469 94236 1555
rect 93796 712 94236 1469
rect 95036 38599 95476 38682
rect 95036 38513 95129 38599
rect 95215 38513 95297 38599
rect 95383 38513 95476 38599
rect 95036 37087 95476 38513
rect 95036 37001 95129 37087
rect 95215 37001 95297 37087
rect 95383 37001 95476 37087
rect 95036 35575 95476 37001
rect 95036 35489 95129 35575
rect 95215 35489 95297 35575
rect 95383 35489 95476 35575
rect 95036 34063 95476 35489
rect 95036 33977 95129 34063
rect 95215 33977 95297 34063
rect 95383 33977 95476 34063
rect 95036 32551 95476 33977
rect 95036 32465 95129 32551
rect 95215 32465 95297 32551
rect 95383 32465 95476 32551
rect 95036 31039 95476 32465
rect 95036 30953 95129 31039
rect 95215 30953 95297 31039
rect 95383 30953 95476 31039
rect 95036 29527 95476 30953
rect 95036 29441 95129 29527
rect 95215 29441 95297 29527
rect 95383 29441 95476 29527
rect 95036 28015 95476 29441
rect 95036 27929 95129 28015
rect 95215 27929 95297 28015
rect 95383 27929 95476 28015
rect 95036 26503 95476 27929
rect 95036 26417 95129 26503
rect 95215 26417 95297 26503
rect 95383 26417 95476 26503
rect 95036 24991 95476 26417
rect 95036 24905 95129 24991
rect 95215 24905 95297 24991
rect 95383 24905 95476 24991
rect 95036 23479 95476 24905
rect 95036 23393 95129 23479
rect 95215 23393 95297 23479
rect 95383 23393 95476 23479
rect 95036 21967 95476 23393
rect 95036 21881 95129 21967
rect 95215 21881 95297 21967
rect 95383 21881 95476 21967
rect 95036 20455 95476 21881
rect 95036 20369 95129 20455
rect 95215 20369 95297 20455
rect 95383 20369 95476 20455
rect 95036 18943 95476 20369
rect 95036 18857 95129 18943
rect 95215 18857 95297 18943
rect 95383 18857 95476 18943
rect 95036 17431 95476 18857
rect 95036 17345 95129 17431
rect 95215 17345 95297 17431
rect 95383 17345 95476 17431
rect 95036 15919 95476 17345
rect 95036 15833 95129 15919
rect 95215 15833 95297 15919
rect 95383 15833 95476 15919
rect 95036 14407 95476 15833
rect 95036 14321 95129 14407
rect 95215 14321 95297 14407
rect 95383 14321 95476 14407
rect 95036 12895 95476 14321
rect 95036 12809 95129 12895
rect 95215 12809 95297 12895
rect 95383 12809 95476 12895
rect 95036 11383 95476 12809
rect 95036 11297 95129 11383
rect 95215 11297 95297 11383
rect 95383 11297 95476 11383
rect 95036 9871 95476 11297
rect 95036 9785 95129 9871
rect 95215 9785 95297 9871
rect 95383 9785 95476 9871
rect 95036 8359 95476 9785
rect 95036 8273 95129 8359
rect 95215 8273 95297 8359
rect 95383 8273 95476 8359
rect 95036 6847 95476 8273
rect 95036 6761 95129 6847
rect 95215 6761 95297 6847
rect 95383 6761 95476 6847
rect 95036 5335 95476 6761
rect 95036 5249 95129 5335
rect 95215 5249 95297 5335
rect 95383 5249 95476 5335
rect 95036 3823 95476 5249
rect 95036 3737 95129 3823
rect 95215 3737 95297 3823
rect 95383 3737 95476 3823
rect 95036 2311 95476 3737
rect 95036 2225 95129 2311
rect 95215 2225 95297 2311
rect 95383 2225 95476 2311
rect 95036 799 95476 2225
rect 95036 713 95129 799
rect 95215 713 95297 799
rect 95383 713 95476 799
rect 95036 630 95476 713
use sg13g2_inv_1  _055_
timestamp 1676382929
transform 1 0 21696 0 1 17388
box -48 -56 336 834
use sg13g2_inv_1  _056_
timestamp 1676382929
transform 1 0 21216 0 1 17388
box -48 -56 336 834
use sg13g2_inv_4  _057_
timestamp 1676383058
transform 1 0 18720 0 1 18900
box -48 -56 624 834
use sg13g2_inv_1  _058_
timestamp 1676382929
transform -1 0 29088 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _059_
timestamp 1676382929
transform -1 0 29376 0 1 21924
box -48 -56 336 834
use sg13g2_inv_1  _060_
timestamp 1676382929
transform -1 0 27552 0 -1 18900
box -48 -56 336 834
use sg13g2_and2_1  _061_
timestamp 1676901763
transform -1 0 28608 0 1 24948
box -48 -56 528 834
use sg13g2_or2_1  _062_
timestamp 1684236171
transform 1 0 19776 0 1 26460
box -48 -56 528 834
use sg13g2_and2_1  _063_
timestamp 1676901763
transform 1 0 19968 0 -1 27972
box -48 -56 528 834
use sg13g2_o21ai_1  _064_
timestamp 1685175443
transform -1 0 20736 0 1 26460
box -48 -56 538 834
use sg13g2_nand2_2  _065_
timestamp 1685180049
transform -1 0 22656 0 -1 18900
box -48 -56 624 834
use sg13g2_nor2_2  _066_
timestamp 1683979924
transform 1 0 19296 0 1 18900
box -48 -56 624 834
use sg13g2_nand3b_1  _067_
timestamp 1676573470
transform -1 0 19776 0 1 20412
box -48 -56 720 834
use sg13g2_nor2b_2  _068_
timestamp 1685188981
transform 1 0 29568 0 -1 24948
box -54 -56 720 834
use sg13g2_a22oi_1  _069_
timestamp 1685173987
transform -1 0 27744 0 -1 30996
box -48 -56 624 834
use sg13g2_inv_4  _070_
timestamp 1676383058
transform 1 0 27360 0 -1 32508
box -48 -56 624 834
use sg13g2_a22oi_1  _071_
timestamp 1685173987
transform 1 0 35520 0 -1 29484
box -48 -56 624 834
use sg13g2_inv_4  _072_
timestamp 1676383058
transform 1 0 36384 0 1 29484
box -48 -56 624 834
use sg13g2_a22oi_1  _073_
timestamp 1685173987
transform 1 0 18048 0 -1 27972
box -48 -56 624 834
use sg13g2_inv_2  _074_
timestamp 1676382947
transform 1 0 18624 0 -1 27972
box -48 -56 432 834
use sg13g2_and2_1  _075_
timestamp 1676901763
transform -1 0 33408 0 1 12852
box -48 -56 528 834
use sg13g2_xor2_1  _076_
timestamp 1677577977
transform -1 0 16032 0 -1 20412
box -48 -56 816 834
use sg13g2_and2_1  _077_
timestamp 1676901763
transform 1 0 18144 0 -1 15876
box -48 -56 528 834
use sg13g2_nor2b_2  _078_
timestamp 1685188981
transform -1 0 29760 0 1 20412
box -54 -56 720 834
use sg13g2_a22oi_1  _079_
timestamp 1685173987
transform 1 0 33696 0 1 15876
box -48 -56 624 834
use sg13g2_o21ai_1  _080_
timestamp 1685175443
transform 1 0 28608 0 1 21924
box -48 -56 538 834
use sg13g2_nor3_1  _081_
timestamp 1676639442
transform 1 0 30240 0 1 20412
box -48 -56 528 834
use sg13g2_a21oi_2  _082_
timestamp 1685174172
transform -1 0 31488 0 1 20412
box -48 -56 816 834
use sg13g2_nand2_1  _083_
timestamp 1676557249
transform 1 0 35136 0 1 21924
box -48 -56 432 834
use sg13g2_nand2_1  _084_
timestamp 1676557249
transform 1 0 34752 0 -1 20412
box -48 -56 432 834
use sg13g2_nand3_1  _085_
timestamp 1683988354
transform 1 0 28512 0 -1 23436
box -48 -56 528 834
use sg13g2_nand2_1  _086_
timestamp 1676557249
transform -1 0 32736 0 1 21924
box -48 -56 432 834
use sg13g2_nand4_1  _087_
timestamp 1685201930
transform 1 0 33984 0 1 21924
box -48 -56 624 834
use sg13g2_nand2_1  _088_
timestamp 1676557249
transform 1 0 35520 0 1 21924
box -48 -56 432 834
use sg13g2_nand4_1  _089_
timestamp 1685201930
transform -1 0 35136 0 1 21924
box -48 -56 624 834
use sg13g2_nand2_1  _090_
timestamp 1676557249
transform 1 0 33600 0 1 17388
box -48 -56 432 834
use sg13g2_nand2_2  _091_
timestamp 1685180049
transform -1 0 34464 0 -1 17388
box -48 -56 624 834
use sg13g2_a22oi_1  _092_
timestamp 1685173987
transform 1 0 27840 0 -1 15876
box -48 -56 624 834
use sg13g2_nand2_1  _093_
timestamp 1676557249
transform -1 0 27072 0 -1 12852
box -48 -56 432 834
use sg13g2_nand2_2  _094_
timestamp 1685180049
transform 1 0 27648 0 -1 12852
box -48 -56 624 834
use sg13g2_nand2_1  _095_
timestamp 1676557249
transform -1 0 26688 0 -1 12852
box -48 -56 432 834
use sg13g2_nand2_2  _096_
timestamp 1685180049
transform 1 0 27072 0 -1 12852
box -48 -56 624 834
use sg13g2_nor2_1  _097_
timestamp 1676627187
transform 1 0 22080 0 1 17388
box -48 -56 432 834
use sg13g2_nand2b_1  _098_
timestamp 1676567195
transform 1 0 21696 0 -1 20412
box -48 -56 528 834
use sg13g2_xor2_1  _099_
timestamp 1677577977
transform -1 0 18144 0 -1 18900
box -48 -56 816 834
use sg13g2_xnor2_1  _100_
timestamp 1677516600
transform -1 0 16512 0 1 17388
box -48 -56 816 834
use sg13g2_nor2_1  _101_
timestamp 1676627187
transform 1 0 15744 0 -1 17388
box -48 -56 432 834
use sg13g2_nand3_1  _102_
timestamp 1683988354
transform 1 0 21024 0 -1 20412
box -48 -56 528 834
use sg13g2_o21ai_1  _103_
timestamp 1685175443
transform 1 0 23040 0 1 20412
box -48 -56 538 834
use sg13g2_o21ai_1  _104_
timestamp 1685175443
transform 1 0 22560 0 1 20412
box -48 -56 538 834
use sg13g2_nor3_1  _105_
timestamp 1676639442
transform 1 0 22464 0 1 17388
box -48 -56 528 834
use sg13g2_nor3_1  _106_
timestamp 1676639442
transform 1 0 21984 0 -1 17388
box -48 -56 528 834
use sg13g2_and2_1  _107_
timestamp 1676901763
transform 1 0 26784 0 -1 27972
box -48 -56 528 834
use sg13g2_inv_1  _108_
timestamp 1676382929
transform 1 0 31104 0 -1 29484
box -48 -56 336 834
use sg13g2_or2_1  _109_
timestamp 1684236171
transform -1 0 30336 0 1 26460
box -48 -56 528 834
use sg13g2_nand3_1  _110_
timestamp 1683988354
transform -1 0 29856 0 1 27972
box -48 -56 528 834
use sg13g2_or2_1  _111_
timestamp 1684236171
transform -1 0 29856 0 1 26460
box -48 -56 528 834
use sg13g2_a21o_1  _112_
timestamp 1677175127
transform 1 0 28704 0 1 27972
box -48 -56 720 834
use sg13g2_nor2b_1  _113_
timestamp 1685181386
transform 1 0 26304 0 -1 27972
box -54 -56 528 834
use sg13g2_a22oi_1  _114_
timestamp 1685173987
transform 1 0 28032 0 1 27972
box -48 -56 624 834
use sg13g2_nor4_1  _115_
timestamp 1676643125
transform -1 0 29760 0 -1 27972
box -48 -56 624 834
use sg13g2_nor4_1  _116_
timestamp 1676643125
transform -1 0 28512 0 -1 26460
box -48 -56 624 834
use sg13g2_and2_1  _117_
timestamp 1676901763
transform -1 0 23616 0 1 27972
box -48 -56 528 834
use sg13g2_nor3_1  _118_
timestamp 1676639442
transform 1 0 21408 0 -1 26460
box -48 -56 528 834
use sg13g2_a21o_1  _119_
timestamp 1677175127
transform 1 0 21984 0 1 27972
box -48 -56 720 834
use sg13g2_and2_1  _120_
timestamp 1676901763
transform 1 0 23232 0 -1 27972
box -48 -56 528 834
use sg13g2_nand2b_1  _121_
timestamp 1676567195
transform -1 0 37440 0 1 15876
box -48 -56 528 834
use sg13g2_mux2_1  _122_
timestamp 1677247768
transform 1 0 36672 0 1 18900
box -48 -56 1008 834
use sg13g2_a22oi_1  _123_
timestamp 1685173987
transform 1 0 26016 0 -1 18900
box -48 -56 624 834
use sg13g2_dfrbpq_1  _124_
timestamp 1746535128
transform 1 0 17664 0 -1 12852
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _125_
timestamp 1746535128
transform 1 0 22464 0 1 11340
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _126_
timestamp 1746535128
transform 1 0 31296 0 -1 17388
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _127_
timestamp 1746535128
transform 1 0 22560 0 1 14364
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _128_
timestamp 1746535128
transform 1 0 15360 0 -1 15876
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _129_
timestamp 1746535128
transform 1 0 24096 0 1 21924
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _130_
timestamp 1746535128
transform 1 0 33984 0 -1 23436
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _131_
timestamp 1746535128
transform 1 0 14880 0 1 21924
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _132_
timestamp 1746535128
transform 1 0 39072 0 1 21924
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _133_
timestamp 1746535128
transform 1 0 37536 0 -1 15876
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _134_
timestamp 1746535128
transform 1 0 38688 0 1 18900
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _135_
timestamp 1746535128
transform -1 0 29280 0 1 30996
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _136_
timestamp 1746535128
transform 1 0 32640 0 -1 30996
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _137_
timestamp 1746535128
transform 1 0 14784 0 -1 26460
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _138_
timestamp 1746535128
transform 1 0 21312 0 1 30996
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _139_
timestamp 1746535128
transform 1 0 34848 0 1 26460
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _140_
timestamp 1746535128
transform 1 0 15264 0 -1 29484
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _141_
timestamp 1746535128
transform 1 0 26688 0 1 17388
box -48 -56 2640 834
use sg13g2_dfrbpq_2  _142_
timestamp 1746535184
transform 1 0 30816 0 -1 12852
box -48 -56 2736 834
use sg13g2_tiehi  _142__32
timestamp 1680000651
transform 1 0 30432 0 -1 12852
box -48 -56 432 834
use sg13g2_dfrbpq_1  _143_
timestamp 1746535128
transform 1 0 19296 0 -1 23436
box -48 -56 2640 834
use sg13g2_buf_1  _157_
timestamp 1676381911
transform -1 0 19008 0 -1 15876
box -48 -56 432 834
use sg13g2_buf_8  clkbuf_0_clk
timestamp 1676451365
transform 1 0 28224 0 -1 21924
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_2_0__f_clk
timestamp 1676451365
transform -1 0 24384 0 -1 20412
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_2_1__f_clk
timestamp 1676451365
transform -1 0 24192 0 -1 24948
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_2_2__f_clk
timestamp 1676451365
transform 1 0 33024 0 1 18900
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_2_3__f_clk
timestamp 1676451365
transform 1 0 33120 0 1 23436
box -48 -56 1296 834
use sg13g2_buf_1  clkload0
timestamp 1676381911
transform 1 0 22752 0 -1 20412
box -48 -56 432 834
use sg13g2_buf_1  clkload1
timestamp 1676381911
transform 1 0 22560 0 -1 24948
box -48 -56 432 834
use sg13g2_buf_1  clkload2
timestamp 1676381911
transform 1 0 32736 0 1 23436
box -48 -56 432 834
use sg13g2_buf_8  fanout11
timestamp 1676451365
transform 1 0 26112 0 -1 26460
box -48 -56 1296 834
use sg13g2_buf_1  fanout12
timestamp 1676381911
transform -1 0 26112 0 -1 26460
box -48 -56 432 834
use sg13g2_buf_8  fanout13
timestamp 1676451365
transform -1 0 39072 0 1 17388
box -48 -56 1296 834
use sg13g2_buf_8  fanout14
timestamp 1676451365
transform -1 0 35520 0 -1 26460
box -48 -56 1296 834
use sg13g2_buf_8  fanout15
timestamp 1676451365
transform 1 0 39456 0 -1 26460
box -48 -56 1296 834
use sg13g2_decap_8  FILLER_0_0
timestamp 1679581782
transform 1 0 576 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_7
timestamp 1679581782
transform 1 0 1248 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_14
timestamp 1679581782
transform 1 0 1920 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_21
timestamp 1679581782
transform 1 0 2592 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_28
timestamp 1679581782
transform 1 0 3264 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_35
timestamp 1679581782
transform 1 0 3936 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_42
timestamp 1679581782
transform 1 0 4608 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_49
timestamp 1679581782
transform 1 0 5280 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_56
timestamp 1679581782
transform 1 0 5952 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_63
timestamp 1679581782
transform 1 0 6624 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_70
timestamp 1679581782
transform 1 0 7296 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_77
timestamp 1679581782
transform 1 0 7968 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_84
timestamp 1679581782
transform 1 0 8640 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_91
timestamp 1679581782
transform 1 0 9312 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_98
timestamp 1679581782
transform 1 0 9984 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_105
timestamp 1679581782
transform 1 0 10656 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_112
timestamp 1679581782
transform 1 0 11328 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_119
timestamp 1679581782
transform 1 0 12000 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_126
timestamp 1679581782
transform 1 0 12672 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_133
timestamp 1679581782
transform 1 0 13344 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_140
timestamp 1679581782
transform 1 0 14016 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_147
timestamp 1679581782
transform 1 0 14688 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_154
timestamp 1679581782
transform 1 0 15360 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_161
timestamp 1679581782
transform 1 0 16032 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_168
timestamp 1679581782
transform 1 0 16704 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_175
timestamp 1679581782
transform 1 0 17376 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_182
timestamp 1679581782
transform 1 0 18048 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_189
timestamp 1679581782
transform 1 0 18720 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_196
timestamp 1679581782
transform 1 0 19392 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_203
timestamp 1679581782
transform 1 0 20064 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_210
timestamp 1679581782
transform 1 0 20736 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_217
timestamp 1679581782
transform 1 0 21408 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_224
timestamp 1679581782
transform 1 0 22080 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_231
timestamp 1679581782
transform 1 0 22752 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_238
timestamp 1679581782
transform 1 0 23424 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_245
timestamp 1679581782
transform 1 0 24096 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_252
timestamp 1679581782
transform 1 0 24768 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_259
timestamp 1679581782
transform 1 0 25440 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_266
timestamp 1679581782
transform 1 0 26112 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_273
timestamp 1679581782
transform 1 0 26784 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_280
timestamp 1679581782
transform 1 0 27456 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_287
timestamp 1679581782
transform 1 0 28128 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_294
timestamp 1679581782
transform 1 0 28800 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_301
timestamp 1679581782
transform 1 0 29472 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_308
timestamp 1679581782
transform 1 0 30144 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_315
timestamp 1679581782
transform 1 0 30816 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_322
timestamp 1679581782
transform 1 0 31488 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_329
timestamp 1679581782
transform 1 0 32160 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_336
timestamp 1679581782
transform 1 0 32832 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_343
timestamp 1679581782
transform 1 0 33504 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_350
timestamp 1679581782
transform 1 0 34176 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_357
timestamp 1679581782
transform 1 0 34848 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_364
timestamp 1679581782
transform 1 0 35520 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_371
timestamp 1679581782
transform 1 0 36192 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_378
timestamp 1679581782
transform 1 0 36864 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_385
timestamp 1679581782
transform 1 0 37536 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_392
timestamp 1679581782
transform 1 0 38208 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_399
timestamp 1679581782
transform 1 0 38880 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_406
timestamp 1679581782
transform 1 0 39552 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_413
timestamp 1679581782
transform 1 0 40224 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_420
timestamp 1679581782
transform 1 0 40896 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_427
timestamp 1679581782
transform 1 0 41568 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_434
timestamp 1679581782
transform 1 0 42240 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_441
timestamp 1679581782
transform 1 0 42912 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_448
timestamp 1679581782
transform 1 0 43584 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_455
timestamp 1679581782
transform 1 0 44256 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_462
timestamp 1679581782
transform 1 0 44928 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_469
timestamp 1679581782
transform 1 0 45600 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_476
timestamp 1679581782
transform 1 0 46272 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_483
timestamp 1679581782
transform 1 0 46944 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_490
timestamp 1679581782
transform 1 0 47616 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_497
timestamp 1679581782
transform 1 0 48288 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_504
timestamp 1679581782
transform 1 0 48960 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_511
timestamp 1679581782
transform 1 0 49632 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_518
timestamp 1679581782
transform 1 0 50304 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_525
timestamp 1679581782
transform 1 0 50976 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_532
timestamp 1679581782
transform 1 0 51648 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_539
timestamp 1679581782
transform 1 0 52320 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_546
timestamp 1679581782
transform 1 0 52992 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_553
timestamp 1679581782
transform 1 0 53664 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_560
timestamp 1679581782
transform 1 0 54336 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_567
timestamp 1679581782
transform 1 0 55008 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_574
timestamp 1679581782
transform 1 0 55680 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_581
timestamp 1679581782
transform 1 0 56352 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_588
timestamp 1679581782
transform 1 0 57024 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_595
timestamp 1679581782
transform 1 0 57696 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_602
timestamp 1679581782
transform 1 0 58368 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_609
timestamp 1679581782
transform 1 0 59040 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_616
timestamp 1679581782
transform 1 0 59712 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_623
timestamp 1679581782
transform 1 0 60384 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_630
timestamp 1679581782
transform 1 0 61056 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_637
timestamp 1679581782
transform 1 0 61728 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_644
timestamp 1679581782
transform 1 0 62400 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_651
timestamp 1679581782
transform 1 0 63072 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_658
timestamp 1679581782
transform 1 0 63744 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_665
timestamp 1679581782
transform 1 0 64416 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_672
timestamp 1679581782
transform 1 0 65088 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_679
timestamp 1679581782
transform 1 0 65760 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_686
timestamp 1679581782
transform 1 0 66432 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_693
timestamp 1679581782
transform 1 0 67104 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_700
timestamp 1679581782
transform 1 0 67776 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_707
timestamp 1679581782
transform 1 0 68448 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_714
timestamp 1679581782
transform 1 0 69120 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_721
timestamp 1679581782
transform 1 0 69792 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_728
timestamp 1679581782
transform 1 0 70464 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_735
timestamp 1679581782
transform 1 0 71136 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_742
timestamp 1679581782
transform 1 0 71808 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_749
timestamp 1679581782
transform 1 0 72480 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_756
timestamp 1679581782
transform 1 0 73152 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_763
timestamp 1679581782
transform 1 0 73824 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_770
timestamp 1679581782
transform 1 0 74496 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_777
timestamp 1679581782
transform 1 0 75168 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_784
timestamp 1679581782
transform 1 0 75840 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_791
timestamp 1679581782
transform 1 0 76512 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_798
timestamp 1679581782
transform 1 0 77184 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_805
timestamp 1679581782
transform 1 0 77856 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_812
timestamp 1679581782
transform 1 0 78528 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_819
timestamp 1679581782
transform 1 0 79200 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_826
timestamp 1679581782
transform 1 0 79872 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_833
timestamp 1679581782
transform 1 0 80544 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_840
timestamp 1679581782
transform 1 0 81216 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_847
timestamp 1679581782
transform 1 0 81888 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_854
timestamp 1679581782
transform 1 0 82560 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_861
timestamp 1679581782
transform 1 0 83232 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_868
timestamp 1679581782
transform 1 0 83904 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_875
timestamp 1679581782
transform 1 0 84576 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_882
timestamp 1679581782
transform 1 0 85248 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_889
timestamp 1679581782
transform 1 0 85920 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_896
timestamp 1679581782
transform 1 0 86592 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_903
timestamp 1679581782
transform 1 0 87264 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_910
timestamp 1679581782
transform 1 0 87936 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_917
timestamp 1679581782
transform 1 0 88608 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_924
timestamp 1679581782
transform 1 0 89280 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_931
timestamp 1679581782
transform 1 0 89952 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_938
timestamp 1679581782
transform 1 0 90624 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_945
timestamp 1679581782
transform 1 0 91296 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_952
timestamp 1679581782
transform 1 0 91968 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_959
timestamp 1679581782
transform 1 0 92640 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_966
timestamp 1679581782
transform 1 0 93312 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_973
timestamp 1679581782
transform 1 0 93984 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_980
timestamp 1679581782
transform 1 0 94656 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_987
timestamp 1679581782
transform 1 0 95328 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_994
timestamp 1679581782
transform 1 0 96000 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_1001
timestamp 1679581782
transform 1 0 96672 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_1008
timestamp 1679581782
transform 1 0 97344 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_1015
timestamp 1679581782
transform 1 0 98016 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_1022
timestamp 1679581782
transform 1 0 98688 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_0
timestamp 1679581782
transform 1 0 576 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_7
timestamp 1679581782
transform 1 0 1248 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_14
timestamp 1679581782
transform 1 0 1920 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_21
timestamp 1679581782
transform 1 0 2592 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_28
timestamp 1679581782
transform 1 0 3264 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_35
timestamp 1679581782
transform 1 0 3936 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_42
timestamp 1679581782
transform 1 0 4608 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_49
timestamp 1679581782
transform 1 0 5280 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_56
timestamp 1679581782
transform 1 0 5952 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_63
timestamp 1679581782
transform 1 0 6624 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_70
timestamp 1679581782
transform 1 0 7296 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_77
timestamp 1679581782
transform 1 0 7968 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_84
timestamp 1679581782
transform 1 0 8640 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_91
timestamp 1679581782
transform 1 0 9312 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_98
timestamp 1679581782
transform 1 0 9984 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_105
timestamp 1679581782
transform 1 0 10656 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_112
timestamp 1679581782
transform 1 0 11328 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_119
timestamp 1679581782
transform 1 0 12000 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_126
timestamp 1679581782
transform 1 0 12672 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_133
timestamp 1679581782
transform 1 0 13344 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_140
timestamp 1679581782
transform 1 0 14016 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_147
timestamp 1679581782
transform 1 0 14688 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_154
timestamp 1679581782
transform 1 0 15360 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_161
timestamp 1679581782
transform 1 0 16032 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_168
timestamp 1679581782
transform 1 0 16704 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_175
timestamp 1679581782
transform 1 0 17376 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_182
timestamp 1679581782
transform 1 0 18048 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_189
timestamp 1679581782
transform 1 0 18720 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_196
timestamp 1679581782
transform 1 0 19392 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_203
timestamp 1679581782
transform 1 0 20064 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_210
timestamp 1679581782
transform 1 0 20736 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_217
timestamp 1679581782
transform 1 0 21408 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_224
timestamp 1679581782
transform 1 0 22080 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_231
timestamp 1679581782
transform 1 0 22752 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_238
timestamp 1679581782
transform 1 0 23424 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_245
timestamp 1679581782
transform 1 0 24096 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_252
timestamp 1679581782
transform 1 0 24768 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_259
timestamp 1679581782
transform 1 0 25440 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_266
timestamp 1679581782
transform 1 0 26112 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_273
timestamp 1679581782
transform 1 0 26784 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_280
timestamp 1679581782
transform 1 0 27456 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_287
timestamp 1679581782
transform 1 0 28128 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_294
timestamp 1679581782
transform 1 0 28800 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_301
timestamp 1679581782
transform 1 0 29472 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_308
timestamp 1679581782
transform 1 0 30144 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_315
timestamp 1679581782
transform 1 0 30816 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_322
timestamp 1679581782
transform 1 0 31488 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_329
timestamp 1679581782
transform 1 0 32160 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_336
timestamp 1679581782
transform 1 0 32832 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_343
timestamp 1679581782
transform 1 0 33504 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_350
timestamp 1679581782
transform 1 0 34176 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_357
timestamp 1679581782
transform 1 0 34848 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_364
timestamp 1679581782
transform 1 0 35520 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_371
timestamp 1679581782
transform 1 0 36192 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_378
timestamp 1679581782
transform 1 0 36864 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_385
timestamp 1679581782
transform 1 0 37536 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_392
timestamp 1679581782
transform 1 0 38208 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_399
timestamp 1679581782
transform 1 0 38880 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_406
timestamp 1679581782
transform 1 0 39552 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_413
timestamp 1679581782
transform 1 0 40224 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_420
timestamp 1679581782
transform 1 0 40896 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_427
timestamp 1679581782
transform 1 0 41568 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_434
timestamp 1679581782
transform 1 0 42240 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_441
timestamp 1679581782
transform 1 0 42912 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_448
timestamp 1679581782
transform 1 0 43584 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_455
timestamp 1679581782
transform 1 0 44256 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_462
timestamp 1679581782
transform 1 0 44928 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_469
timestamp 1679581782
transform 1 0 45600 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_476
timestamp 1679581782
transform 1 0 46272 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_483
timestamp 1679581782
transform 1 0 46944 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_490
timestamp 1679581782
transform 1 0 47616 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_497
timestamp 1679581782
transform 1 0 48288 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_504
timestamp 1679581782
transform 1 0 48960 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_511
timestamp 1679581782
transform 1 0 49632 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_518
timestamp 1679581782
transform 1 0 50304 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_525
timestamp 1679581782
transform 1 0 50976 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_532
timestamp 1679581782
transform 1 0 51648 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_539
timestamp 1679581782
transform 1 0 52320 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_546
timestamp 1679581782
transform 1 0 52992 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_553
timestamp 1679581782
transform 1 0 53664 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_560
timestamp 1679581782
transform 1 0 54336 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_567
timestamp 1679581782
transform 1 0 55008 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_574
timestamp 1679581782
transform 1 0 55680 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_581
timestamp 1679581782
transform 1 0 56352 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_588
timestamp 1679581782
transform 1 0 57024 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_595
timestamp 1679581782
transform 1 0 57696 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_602
timestamp 1679581782
transform 1 0 58368 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_609
timestamp 1679581782
transform 1 0 59040 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_616
timestamp 1679581782
transform 1 0 59712 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_623
timestamp 1679581782
transform 1 0 60384 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_630
timestamp 1679581782
transform 1 0 61056 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_637
timestamp 1679581782
transform 1 0 61728 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_644
timestamp 1679581782
transform 1 0 62400 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_651
timestamp 1679581782
transform 1 0 63072 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_658
timestamp 1679581782
transform 1 0 63744 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_665
timestamp 1679581782
transform 1 0 64416 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_672
timestamp 1679581782
transform 1 0 65088 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_679
timestamp 1679581782
transform 1 0 65760 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_686
timestamp 1679581782
transform 1 0 66432 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_693
timestamp 1679581782
transform 1 0 67104 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_700
timestamp 1679581782
transform 1 0 67776 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_707
timestamp 1679581782
transform 1 0 68448 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_714
timestamp 1679581782
transform 1 0 69120 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_721
timestamp 1679581782
transform 1 0 69792 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_728
timestamp 1679581782
transform 1 0 70464 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_735
timestamp 1679581782
transform 1 0 71136 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_742
timestamp 1679581782
transform 1 0 71808 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_749
timestamp 1679581782
transform 1 0 72480 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_756
timestamp 1679581782
transform 1 0 73152 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_763
timestamp 1679581782
transform 1 0 73824 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_770
timestamp 1679581782
transform 1 0 74496 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_777
timestamp 1679581782
transform 1 0 75168 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_784
timestamp 1679581782
transform 1 0 75840 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_791
timestamp 1679581782
transform 1 0 76512 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_798
timestamp 1679581782
transform 1 0 77184 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_805
timestamp 1679581782
transform 1 0 77856 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_812
timestamp 1679581782
transform 1 0 78528 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_819
timestamp 1679581782
transform 1 0 79200 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_826
timestamp 1679581782
transform 1 0 79872 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_833
timestamp 1679581782
transform 1 0 80544 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_840
timestamp 1679581782
transform 1 0 81216 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_847
timestamp 1679581782
transform 1 0 81888 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_854
timestamp 1679581782
transform 1 0 82560 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_861
timestamp 1679581782
transform 1 0 83232 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_868
timestamp 1679581782
transform 1 0 83904 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_875
timestamp 1679581782
transform 1 0 84576 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_882
timestamp 1679581782
transform 1 0 85248 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_889
timestamp 1679581782
transform 1 0 85920 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_896
timestamp 1679581782
transform 1 0 86592 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_903
timestamp 1679581782
transform 1 0 87264 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_910
timestamp 1679581782
transform 1 0 87936 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_917
timestamp 1679581782
transform 1 0 88608 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_924
timestamp 1679581782
transform 1 0 89280 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_931
timestamp 1679581782
transform 1 0 89952 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_938
timestamp 1679581782
transform 1 0 90624 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_945
timestamp 1679581782
transform 1 0 91296 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_952
timestamp 1679581782
transform 1 0 91968 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_959
timestamp 1679581782
transform 1 0 92640 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_966
timestamp 1679581782
transform 1 0 93312 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_973
timestamp 1679581782
transform 1 0 93984 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_980
timestamp 1679581782
transform 1 0 94656 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_987
timestamp 1679581782
transform 1 0 95328 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_994
timestamp 1679581782
transform 1 0 96000 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_1001
timestamp 1679581782
transform 1 0 96672 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_1008
timestamp 1679581782
transform 1 0 97344 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_1015
timestamp 1679581782
transform 1 0 98016 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_1022
timestamp 1679581782
transform 1 0 98688 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_4
timestamp 1679581782
transform 1 0 960 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_11
timestamp 1679581782
transform 1 0 1632 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_18
timestamp 1679581782
transform 1 0 2304 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_25
timestamp 1679581782
transform 1 0 2976 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_32
timestamp 1679581782
transform 1 0 3648 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_39
timestamp 1679581782
transform 1 0 4320 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_46
timestamp 1679581782
transform 1 0 4992 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_53
timestamp 1679581782
transform 1 0 5664 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_60
timestamp 1679581782
transform 1 0 6336 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_67
timestamp 1679581782
transform 1 0 7008 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_74
timestamp 1679581782
transform 1 0 7680 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_81
timestamp 1679581782
transform 1 0 8352 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_88
timestamp 1679581782
transform 1 0 9024 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_95
timestamp 1679581782
transform 1 0 9696 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_102
timestamp 1679581782
transform 1 0 10368 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_109
timestamp 1679581782
transform 1 0 11040 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_116
timestamp 1679581782
transform 1 0 11712 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_123
timestamp 1679581782
transform 1 0 12384 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_130
timestamp 1679581782
transform 1 0 13056 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_137
timestamp 1679581782
transform 1 0 13728 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_144
timestamp 1679581782
transform 1 0 14400 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_151
timestamp 1679581782
transform 1 0 15072 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_158
timestamp 1679581782
transform 1 0 15744 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_165
timestamp 1679581782
transform 1 0 16416 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_172
timestamp 1679581782
transform 1 0 17088 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_179
timestamp 1679581782
transform 1 0 17760 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_186
timestamp 1679581782
transform 1 0 18432 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_193
timestamp 1679581782
transform 1 0 19104 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_200
timestamp 1679581782
transform 1 0 19776 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_207
timestamp 1679581782
transform 1 0 20448 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_214
timestamp 1679581782
transform 1 0 21120 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_221
timestamp 1679581782
transform 1 0 21792 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_228
timestamp 1679581782
transform 1 0 22464 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_235
timestamp 1679581782
transform 1 0 23136 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_242
timestamp 1679581782
transform 1 0 23808 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_249
timestamp 1679581782
transform 1 0 24480 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_256
timestamp 1679581782
transform 1 0 25152 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_263
timestamp 1679581782
transform 1 0 25824 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_270
timestamp 1679581782
transform 1 0 26496 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_277
timestamp 1679581782
transform 1 0 27168 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_284
timestamp 1679581782
transform 1 0 27840 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_291
timestamp 1679581782
transform 1 0 28512 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_298
timestamp 1679581782
transform 1 0 29184 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_305
timestamp 1679581782
transform 1 0 29856 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_312
timestamp 1679581782
transform 1 0 30528 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_319
timestamp 1679581782
transform 1 0 31200 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_326
timestamp 1679581782
transform 1 0 31872 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_333
timestamp 1679581782
transform 1 0 32544 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_340
timestamp 1679581782
transform 1 0 33216 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_347
timestamp 1679581782
transform 1 0 33888 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_354
timestamp 1679581782
transform 1 0 34560 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_361
timestamp 1679581782
transform 1 0 35232 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_368
timestamp 1679581782
transform 1 0 35904 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_375
timestamp 1679581782
transform 1 0 36576 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_382
timestamp 1679581782
transform 1 0 37248 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_389
timestamp 1679581782
transform 1 0 37920 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_396
timestamp 1679581782
transform 1 0 38592 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_403
timestamp 1679581782
transform 1 0 39264 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_410
timestamp 1679581782
transform 1 0 39936 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_417
timestamp 1679581782
transform 1 0 40608 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_424
timestamp 1679581782
transform 1 0 41280 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_431
timestamp 1679581782
transform 1 0 41952 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_438
timestamp 1679581782
transform 1 0 42624 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_445
timestamp 1679581782
transform 1 0 43296 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_452
timestamp 1679581782
transform 1 0 43968 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_459
timestamp 1679581782
transform 1 0 44640 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_466
timestamp 1679581782
transform 1 0 45312 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_473
timestamp 1679581782
transform 1 0 45984 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_480
timestamp 1679581782
transform 1 0 46656 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_487
timestamp 1679581782
transform 1 0 47328 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_494
timestamp 1679581782
transform 1 0 48000 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_501
timestamp 1679581782
transform 1 0 48672 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_508
timestamp 1679581782
transform 1 0 49344 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_515
timestamp 1679581782
transform 1 0 50016 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_522
timestamp 1679581782
transform 1 0 50688 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_529
timestamp 1679581782
transform 1 0 51360 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_536
timestamp 1679581782
transform 1 0 52032 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_543
timestamp 1679581782
transform 1 0 52704 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_550
timestamp 1679581782
transform 1 0 53376 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_557
timestamp 1679581782
transform 1 0 54048 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_564
timestamp 1679581782
transform 1 0 54720 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_571
timestamp 1679581782
transform 1 0 55392 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_578
timestamp 1679581782
transform 1 0 56064 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_585
timestamp 1679581782
transform 1 0 56736 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_592
timestamp 1679581782
transform 1 0 57408 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_599
timestamp 1679581782
transform 1 0 58080 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_606
timestamp 1679581782
transform 1 0 58752 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_613
timestamp 1679581782
transform 1 0 59424 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_620
timestamp 1679581782
transform 1 0 60096 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_627
timestamp 1679581782
transform 1 0 60768 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_634
timestamp 1679581782
transform 1 0 61440 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_641
timestamp 1679581782
transform 1 0 62112 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_648
timestamp 1679581782
transform 1 0 62784 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_655
timestamp 1679581782
transform 1 0 63456 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_662
timestamp 1679581782
transform 1 0 64128 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_669
timestamp 1679581782
transform 1 0 64800 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_676
timestamp 1679581782
transform 1 0 65472 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_683
timestamp 1679581782
transform 1 0 66144 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_690
timestamp 1679581782
transform 1 0 66816 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_697
timestamp 1679581782
transform 1 0 67488 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_704
timestamp 1679581782
transform 1 0 68160 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_711
timestamp 1679581782
transform 1 0 68832 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_718
timestamp 1679581782
transform 1 0 69504 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_725
timestamp 1679581782
transform 1 0 70176 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_732
timestamp 1679581782
transform 1 0 70848 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_739
timestamp 1679581782
transform 1 0 71520 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_746
timestamp 1679581782
transform 1 0 72192 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_753
timestamp 1679581782
transform 1 0 72864 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_760
timestamp 1679581782
transform 1 0 73536 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_767
timestamp 1679581782
transform 1 0 74208 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_774
timestamp 1679581782
transform 1 0 74880 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_781
timestamp 1679581782
transform 1 0 75552 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_788
timestamp 1679581782
transform 1 0 76224 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_795
timestamp 1679581782
transform 1 0 76896 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_802
timestamp 1679581782
transform 1 0 77568 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_809
timestamp 1679581782
transform 1 0 78240 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_816
timestamp 1679581782
transform 1 0 78912 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_823
timestamp 1679581782
transform 1 0 79584 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_830
timestamp 1679581782
transform 1 0 80256 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_837
timestamp 1679581782
transform 1 0 80928 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_844
timestamp 1679581782
transform 1 0 81600 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_851
timestamp 1679581782
transform 1 0 82272 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_858
timestamp 1679581782
transform 1 0 82944 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_865
timestamp 1679581782
transform 1 0 83616 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_872
timestamp 1679581782
transform 1 0 84288 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_879
timestamp 1679581782
transform 1 0 84960 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_886
timestamp 1679581782
transform 1 0 85632 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_893
timestamp 1679581782
transform 1 0 86304 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_900
timestamp 1679581782
transform 1 0 86976 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_907
timestamp 1679581782
transform 1 0 87648 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_914
timestamp 1679581782
transform 1 0 88320 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_921
timestamp 1679581782
transform 1 0 88992 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_928
timestamp 1679581782
transform 1 0 89664 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_935
timestamp 1679581782
transform 1 0 90336 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_942
timestamp 1679581782
transform 1 0 91008 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_949
timestamp 1679581782
transform 1 0 91680 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_956
timestamp 1679581782
transform 1 0 92352 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_963
timestamp 1679581782
transform 1 0 93024 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_970
timestamp 1679581782
transform 1 0 93696 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_977
timestamp 1679581782
transform 1 0 94368 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_984
timestamp 1679581782
transform 1 0 95040 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_991
timestamp 1679581782
transform 1 0 95712 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_998
timestamp 1679581782
transform 1 0 96384 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_1005
timestamp 1679581782
transform 1 0 97056 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_1012
timestamp 1679581782
transform 1 0 97728 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_1019
timestamp 1679581782
transform 1 0 98400 0 1 2268
box -48 -56 720 834
use sg13g2_fill_2  FILLER_2_1026
timestamp 1677580104
transform 1 0 99072 0 1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_1028
timestamp 1677579658
transform 1 0 99264 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_4
timestamp 1679581782
transform 1 0 960 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_11
timestamp 1679581782
transform 1 0 1632 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_18
timestamp 1679581782
transform 1 0 2304 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_25
timestamp 1679581782
transform 1 0 2976 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_32
timestamp 1679581782
transform 1 0 3648 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_39
timestamp 1679581782
transform 1 0 4320 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_46
timestamp 1679581782
transform 1 0 4992 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_53
timestamp 1679581782
transform 1 0 5664 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_60
timestamp 1679581782
transform 1 0 6336 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_67
timestamp 1679581782
transform 1 0 7008 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_74
timestamp 1679581782
transform 1 0 7680 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_81
timestamp 1679581782
transform 1 0 8352 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_88
timestamp 1679581782
transform 1 0 9024 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_95
timestamp 1679581782
transform 1 0 9696 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_102
timestamp 1679581782
transform 1 0 10368 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_109
timestamp 1679581782
transform 1 0 11040 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_116
timestamp 1679581782
transform 1 0 11712 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_123
timestamp 1679581782
transform 1 0 12384 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_130
timestamp 1679581782
transform 1 0 13056 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_137
timestamp 1679581782
transform 1 0 13728 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_144
timestamp 1679581782
transform 1 0 14400 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_151
timestamp 1679581782
transform 1 0 15072 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_158
timestamp 1679581782
transform 1 0 15744 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_165
timestamp 1679581782
transform 1 0 16416 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_172
timestamp 1679581782
transform 1 0 17088 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_179
timestamp 1679581782
transform 1 0 17760 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_186
timestamp 1679581782
transform 1 0 18432 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_193
timestamp 1679581782
transform 1 0 19104 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_200
timestamp 1679581782
transform 1 0 19776 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_207
timestamp 1679581782
transform 1 0 20448 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_214
timestamp 1679581782
transform 1 0 21120 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_221
timestamp 1679581782
transform 1 0 21792 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_228
timestamp 1679581782
transform 1 0 22464 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_235
timestamp 1679581782
transform 1 0 23136 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_242
timestamp 1679581782
transform 1 0 23808 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_249
timestamp 1679581782
transform 1 0 24480 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_256
timestamp 1679581782
transform 1 0 25152 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_263
timestamp 1679581782
transform 1 0 25824 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_270
timestamp 1679581782
transform 1 0 26496 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_277
timestamp 1679581782
transform 1 0 27168 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_284
timestamp 1679581782
transform 1 0 27840 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_291
timestamp 1679581782
transform 1 0 28512 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_298
timestamp 1679581782
transform 1 0 29184 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_305
timestamp 1679581782
transform 1 0 29856 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_312
timestamp 1679581782
transform 1 0 30528 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_319
timestamp 1679581782
transform 1 0 31200 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_326
timestamp 1679581782
transform 1 0 31872 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_333
timestamp 1679581782
transform 1 0 32544 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_340
timestamp 1679581782
transform 1 0 33216 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_347
timestamp 1679581782
transform 1 0 33888 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_354
timestamp 1679581782
transform 1 0 34560 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_361
timestamp 1679581782
transform 1 0 35232 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_368
timestamp 1679581782
transform 1 0 35904 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_375
timestamp 1679581782
transform 1 0 36576 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_382
timestamp 1679581782
transform 1 0 37248 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_389
timestamp 1679581782
transform 1 0 37920 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_396
timestamp 1679581782
transform 1 0 38592 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_403
timestamp 1679581782
transform 1 0 39264 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_410
timestamp 1679581782
transform 1 0 39936 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_417
timestamp 1679581782
transform 1 0 40608 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_424
timestamp 1679581782
transform 1 0 41280 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_431
timestamp 1679581782
transform 1 0 41952 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_438
timestamp 1679581782
transform 1 0 42624 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_445
timestamp 1679581782
transform 1 0 43296 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_452
timestamp 1679581782
transform 1 0 43968 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_459
timestamp 1679581782
transform 1 0 44640 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_466
timestamp 1679581782
transform 1 0 45312 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_473
timestamp 1679581782
transform 1 0 45984 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_480
timestamp 1679581782
transform 1 0 46656 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_487
timestamp 1679581782
transform 1 0 47328 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_494
timestamp 1679581782
transform 1 0 48000 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_501
timestamp 1679581782
transform 1 0 48672 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_508
timestamp 1679581782
transform 1 0 49344 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_515
timestamp 1679581782
transform 1 0 50016 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_522
timestamp 1679581782
transform 1 0 50688 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_529
timestamp 1679581782
transform 1 0 51360 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_536
timestamp 1679581782
transform 1 0 52032 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_543
timestamp 1679581782
transform 1 0 52704 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_550
timestamp 1679581782
transform 1 0 53376 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_557
timestamp 1679581782
transform 1 0 54048 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_564
timestamp 1679581782
transform 1 0 54720 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_571
timestamp 1679581782
transform 1 0 55392 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_578
timestamp 1679581782
transform 1 0 56064 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_585
timestamp 1679581782
transform 1 0 56736 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_592
timestamp 1679581782
transform 1 0 57408 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_599
timestamp 1679581782
transform 1 0 58080 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_606
timestamp 1679581782
transform 1 0 58752 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_613
timestamp 1679581782
transform 1 0 59424 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_620
timestamp 1679581782
transform 1 0 60096 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_627
timestamp 1679581782
transform 1 0 60768 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_634
timestamp 1679581782
transform 1 0 61440 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_641
timestamp 1679581782
transform 1 0 62112 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_648
timestamp 1679581782
transform 1 0 62784 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_655
timestamp 1679581782
transform 1 0 63456 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_662
timestamp 1679581782
transform 1 0 64128 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_669
timestamp 1679581782
transform 1 0 64800 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_676
timestamp 1679581782
transform 1 0 65472 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_683
timestamp 1679581782
transform 1 0 66144 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_690
timestamp 1679581782
transform 1 0 66816 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_697
timestamp 1679581782
transform 1 0 67488 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_704
timestamp 1679581782
transform 1 0 68160 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_711
timestamp 1679581782
transform 1 0 68832 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_718
timestamp 1679581782
transform 1 0 69504 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_725
timestamp 1679581782
transform 1 0 70176 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_732
timestamp 1679581782
transform 1 0 70848 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_739
timestamp 1679581782
transform 1 0 71520 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_746
timestamp 1679581782
transform 1 0 72192 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_753
timestamp 1679581782
transform 1 0 72864 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_760
timestamp 1679581782
transform 1 0 73536 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_767
timestamp 1679581782
transform 1 0 74208 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_774
timestamp 1679581782
transform 1 0 74880 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_781
timestamp 1679581782
transform 1 0 75552 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_788
timestamp 1679581782
transform 1 0 76224 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_795
timestamp 1679581782
transform 1 0 76896 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_802
timestamp 1679581782
transform 1 0 77568 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_809
timestamp 1679581782
transform 1 0 78240 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_816
timestamp 1679581782
transform 1 0 78912 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_823
timestamp 1679581782
transform 1 0 79584 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_830
timestamp 1679581782
transform 1 0 80256 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_837
timestamp 1679581782
transform 1 0 80928 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_844
timestamp 1679581782
transform 1 0 81600 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_851
timestamp 1679581782
transform 1 0 82272 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_858
timestamp 1679581782
transform 1 0 82944 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_865
timestamp 1679581782
transform 1 0 83616 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_872
timestamp 1679581782
transform 1 0 84288 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_879
timestamp 1679581782
transform 1 0 84960 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_886
timestamp 1679581782
transform 1 0 85632 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_893
timestamp 1679581782
transform 1 0 86304 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_900
timestamp 1679581782
transform 1 0 86976 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_907
timestamp 1679581782
transform 1 0 87648 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_914
timestamp 1679581782
transform 1 0 88320 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_921
timestamp 1679581782
transform 1 0 88992 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_928
timestamp 1679581782
transform 1 0 89664 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_935
timestamp 1679581782
transform 1 0 90336 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_942
timestamp 1679581782
transform 1 0 91008 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_949
timestamp 1679581782
transform 1 0 91680 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_956
timestamp 1679581782
transform 1 0 92352 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_963
timestamp 1679581782
transform 1 0 93024 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_970
timestamp 1679581782
transform 1 0 93696 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_977
timestamp 1679581782
transform 1 0 94368 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_984
timestamp 1679581782
transform 1 0 95040 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_991
timestamp 1679581782
transform 1 0 95712 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_998
timestamp 1679581782
transform 1 0 96384 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_1005
timestamp 1679581782
transform 1 0 97056 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_1012
timestamp 1679581782
transform 1 0 97728 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_1019
timestamp 1679581782
transform 1 0 98400 0 -1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_3_1026
timestamp 1677580104
transform 1 0 99072 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_1028
timestamp 1677579658
transform 1 0 99264 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_4
timestamp 1679581782
transform 1 0 960 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_11
timestamp 1679581782
transform 1 0 1632 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_18
timestamp 1679581782
transform 1 0 2304 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_25
timestamp 1679581782
transform 1 0 2976 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_32
timestamp 1679581782
transform 1 0 3648 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_39
timestamp 1679581782
transform 1 0 4320 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_46
timestamp 1679581782
transform 1 0 4992 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_53
timestamp 1679581782
transform 1 0 5664 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_60
timestamp 1679581782
transform 1 0 6336 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_67
timestamp 1679581782
transform 1 0 7008 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_74
timestamp 1679581782
transform 1 0 7680 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_81
timestamp 1679581782
transform 1 0 8352 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_88
timestamp 1679581782
transform 1 0 9024 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_95
timestamp 1679581782
transform 1 0 9696 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_102
timestamp 1679581782
transform 1 0 10368 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_109
timestamp 1679581782
transform 1 0 11040 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_116
timestamp 1679581782
transform 1 0 11712 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_123
timestamp 1679581782
transform 1 0 12384 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_130
timestamp 1679581782
transform 1 0 13056 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_137
timestamp 1679581782
transform 1 0 13728 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_144
timestamp 1679581782
transform 1 0 14400 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_151
timestamp 1679581782
transform 1 0 15072 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_158
timestamp 1679581782
transform 1 0 15744 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_165
timestamp 1679581782
transform 1 0 16416 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_172
timestamp 1679581782
transform 1 0 17088 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_179
timestamp 1679581782
transform 1 0 17760 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_186
timestamp 1679581782
transform 1 0 18432 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_193
timestamp 1679581782
transform 1 0 19104 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_200
timestamp 1679581782
transform 1 0 19776 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_207
timestamp 1679581782
transform 1 0 20448 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_214
timestamp 1679581782
transform 1 0 21120 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_221
timestamp 1679581782
transform 1 0 21792 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_228
timestamp 1679581782
transform 1 0 22464 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_235
timestamp 1679581782
transform 1 0 23136 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_242
timestamp 1679581782
transform 1 0 23808 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_249
timestamp 1679581782
transform 1 0 24480 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_256
timestamp 1679581782
transform 1 0 25152 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_263
timestamp 1679581782
transform 1 0 25824 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_270
timestamp 1679581782
transform 1 0 26496 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_277
timestamp 1679581782
transform 1 0 27168 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_284
timestamp 1679581782
transform 1 0 27840 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_291
timestamp 1679581782
transform 1 0 28512 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_298
timestamp 1679581782
transform 1 0 29184 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_305
timestamp 1679581782
transform 1 0 29856 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_312
timestamp 1679581782
transform 1 0 30528 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_319
timestamp 1679581782
transform 1 0 31200 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_326
timestamp 1679581782
transform 1 0 31872 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_333
timestamp 1679581782
transform 1 0 32544 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_340
timestamp 1679581782
transform 1 0 33216 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_347
timestamp 1679581782
transform 1 0 33888 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_354
timestamp 1679581782
transform 1 0 34560 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_361
timestamp 1679581782
transform 1 0 35232 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_368
timestamp 1679581782
transform 1 0 35904 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_375
timestamp 1679581782
transform 1 0 36576 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_382
timestamp 1679581782
transform 1 0 37248 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_389
timestamp 1679581782
transform 1 0 37920 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_396
timestamp 1679581782
transform 1 0 38592 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_403
timestamp 1679581782
transform 1 0 39264 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_410
timestamp 1679581782
transform 1 0 39936 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_417
timestamp 1679581782
transform 1 0 40608 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_424
timestamp 1679581782
transform 1 0 41280 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_431
timestamp 1679581782
transform 1 0 41952 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_438
timestamp 1679581782
transform 1 0 42624 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_445
timestamp 1679581782
transform 1 0 43296 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_452
timestamp 1679581782
transform 1 0 43968 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_459
timestamp 1679581782
transform 1 0 44640 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_466
timestamp 1679581782
transform 1 0 45312 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_473
timestamp 1679581782
transform 1 0 45984 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_480
timestamp 1679581782
transform 1 0 46656 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_487
timestamp 1679581782
transform 1 0 47328 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_494
timestamp 1679581782
transform 1 0 48000 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_501
timestamp 1679581782
transform 1 0 48672 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_508
timestamp 1679581782
transform 1 0 49344 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_515
timestamp 1679581782
transform 1 0 50016 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_522
timestamp 1679581782
transform 1 0 50688 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_529
timestamp 1679581782
transform 1 0 51360 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_536
timestamp 1679581782
transform 1 0 52032 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_543
timestamp 1679581782
transform 1 0 52704 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_550
timestamp 1679581782
transform 1 0 53376 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_557
timestamp 1679581782
transform 1 0 54048 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_564
timestamp 1679581782
transform 1 0 54720 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_571
timestamp 1679581782
transform 1 0 55392 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_578
timestamp 1679581782
transform 1 0 56064 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_585
timestamp 1679581782
transform 1 0 56736 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_592
timestamp 1679581782
transform 1 0 57408 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_599
timestamp 1679581782
transform 1 0 58080 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_606
timestamp 1679581782
transform 1 0 58752 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_613
timestamp 1679581782
transform 1 0 59424 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_620
timestamp 1679581782
transform 1 0 60096 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_627
timestamp 1679581782
transform 1 0 60768 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_634
timestamp 1679581782
transform 1 0 61440 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_641
timestamp 1679581782
transform 1 0 62112 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_648
timestamp 1679581782
transform 1 0 62784 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_655
timestamp 1679581782
transform 1 0 63456 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_662
timestamp 1679581782
transform 1 0 64128 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_669
timestamp 1679581782
transform 1 0 64800 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_676
timestamp 1679581782
transform 1 0 65472 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_683
timestamp 1679581782
transform 1 0 66144 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_690
timestamp 1679581782
transform 1 0 66816 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_697
timestamp 1679581782
transform 1 0 67488 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_704
timestamp 1679581782
transform 1 0 68160 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_711
timestamp 1679581782
transform 1 0 68832 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_718
timestamp 1679581782
transform 1 0 69504 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_725
timestamp 1679581782
transform 1 0 70176 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_732
timestamp 1679581782
transform 1 0 70848 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_739
timestamp 1679581782
transform 1 0 71520 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_746
timestamp 1679581782
transform 1 0 72192 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_753
timestamp 1679581782
transform 1 0 72864 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_760
timestamp 1679581782
transform 1 0 73536 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_767
timestamp 1679581782
transform 1 0 74208 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_774
timestamp 1679581782
transform 1 0 74880 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_781
timestamp 1679581782
transform 1 0 75552 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_788
timestamp 1679581782
transform 1 0 76224 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_795
timestamp 1679581782
transform 1 0 76896 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_802
timestamp 1679581782
transform 1 0 77568 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_809
timestamp 1679581782
transform 1 0 78240 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_816
timestamp 1679581782
transform 1 0 78912 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_823
timestamp 1679581782
transform 1 0 79584 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_830
timestamp 1679581782
transform 1 0 80256 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_837
timestamp 1679581782
transform 1 0 80928 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_844
timestamp 1679581782
transform 1 0 81600 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_851
timestamp 1679581782
transform 1 0 82272 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_858
timestamp 1679581782
transform 1 0 82944 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_865
timestamp 1679581782
transform 1 0 83616 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_872
timestamp 1679581782
transform 1 0 84288 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_879
timestamp 1679581782
transform 1 0 84960 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_886
timestamp 1679581782
transform 1 0 85632 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_893
timestamp 1679581782
transform 1 0 86304 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_900
timestamp 1679581782
transform 1 0 86976 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_907
timestamp 1679581782
transform 1 0 87648 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_914
timestamp 1679581782
transform 1 0 88320 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_921
timestamp 1679581782
transform 1 0 88992 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_928
timestamp 1679581782
transform 1 0 89664 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_935
timestamp 1679581782
transform 1 0 90336 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_942
timestamp 1679581782
transform 1 0 91008 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_949
timestamp 1679581782
transform 1 0 91680 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_956
timestamp 1679581782
transform 1 0 92352 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_963
timestamp 1679581782
transform 1 0 93024 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_970
timestamp 1679581782
transform 1 0 93696 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_977
timestamp 1679581782
transform 1 0 94368 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_984
timestamp 1679581782
transform 1 0 95040 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_991
timestamp 1679581782
transform 1 0 95712 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_998
timestamp 1679581782
transform 1 0 96384 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_1005
timestamp 1679581782
transform 1 0 97056 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_1012
timestamp 1679581782
transform 1 0 97728 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_1019
timestamp 1679581782
transform 1 0 98400 0 1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_4_1026
timestamp 1677580104
transform 1 0 99072 0 1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_1028
timestamp 1677579658
transform 1 0 99264 0 1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_4
timestamp 1679581782
transform 1 0 960 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_11
timestamp 1679581782
transform 1 0 1632 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_18
timestamp 1679581782
transform 1 0 2304 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_25
timestamp 1679581782
transform 1 0 2976 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_32
timestamp 1679581782
transform 1 0 3648 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_39
timestamp 1679581782
transform 1 0 4320 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_46
timestamp 1679581782
transform 1 0 4992 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_53
timestamp 1679581782
transform 1 0 5664 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_60
timestamp 1679581782
transform 1 0 6336 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_67
timestamp 1679581782
transform 1 0 7008 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_74
timestamp 1679581782
transform 1 0 7680 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_81
timestamp 1679581782
transform 1 0 8352 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_88
timestamp 1679581782
transform 1 0 9024 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_95
timestamp 1679581782
transform 1 0 9696 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_102
timestamp 1679581782
transform 1 0 10368 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_109
timestamp 1679581782
transform 1 0 11040 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_116
timestamp 1679581782
transform 1 0 11712 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_123
timestamp 1679581782
transform 1 0 12384 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_130
timestamp 1679581782
transform 1 0 13056 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_137
timestamp 1679581782
transform 1 0 13728 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_144
timestamp 1679581782
transform 1 0 14400 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_151
timestamp 1679581782
transform 1 0 15072 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_158
timestamp 1679581782
transform 1 0 15744 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_165
timestamp 1679581782
transform 1 0 16416 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_172
timestamp 1679581782
transform 1 0 17088 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_179
timestamp 1679581782
transform 1 0 17760 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_186
timestamp 1679581782
transform 1 0 18432 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_193
timestamp 1679581782
transform 1 0 19104 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_200
timestamp 1679581782
transform 1 0 19776 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_207
timestamp 1679581782
transform 1 0 20448 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_214
timestamp 1679581782
transform 1 0 21120 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_221
timestamp 1679581782
transform 1 0 21792 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_228
timestamp 1679581782
transform 1 0 22464 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_235
timestamp 1679581782
transform 1 0 23136 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_242
timestamp 1679581782
transform 1 0 23808 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_249
timestamp 1679581782
transform 1 0 24480 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_256
timestamp 1679581782
transform 1 0 25152 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_263
timestamp 1679581782
transform 1 0 25824 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_270
timestamp 1679581782
transform 1 0 26496 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_277
timestamp 1679581782
transform 1 0 27168 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_284
timestamp 1679581782
transform 1 0 27840 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_291
timestamp 1679581782
transform 1 0 28512 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_298
timestamp 1679581782
transform 1 0 29184 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_305
timestamp 1679581782
transform 1 0 29856 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_312
timestamp 1679581782
transform 1 0 30528 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_319
timestamp 1679581782
transform 1 0 31200 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_326
timestamp 1679581782
transform 1 0 31872 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_333
timestamp 1679581782
transform 1 0 32544 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_340
timestamp 1679581782
transform 1 0 33216 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_347
timestamp 1679581782
transform 1 0 33888 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_354
timestamp 1679581782
transform 1 0 34560 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_361
timestamp 1679581782
transform 1 0 35232 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_368
timestamp 1679581782
transform 1 0 35904 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_375
timestamp 1679581782
transform 1 0 36576 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_382
timestamp 1679581782
transform 1 0 37248 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_389
timestamp 1679581782
transform 1 0 37920 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_396
timestamp 1679581782
transform 1 0 38592 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_403
timestamp 1679581782
transform 1 0 39264 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_410
timestamp 1679581782
transform 1 0 39936 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_417
timestamp 1679581782
transform 1 0 40608 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_424
timestamp 1679581782
transform 1 0 41280 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_431
timestamp 1679581782
transform 1 0 41952 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_438
timestamp 1679581782
transform 1 0 42624 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_445
timestamp 1679581782
transform 1 0 43296 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_452
timestamp 1679581782
transform 1 0 43968 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_459
timestamp 1679581782
transform 1 0 44640 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_466
timestamp 1679581782
transform 1 0 45312 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_473
timestamp 1679581782
transform 1 0 45984 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_480
timestamp 1679581782
transform 1 0 46656 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_487
timestamp 1679581782
transform 1 0 47328 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_494
timestamp 1679581782
transform 1 0 48000 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_501
timestamp 1679581782
transform 1 0 48672 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_508
timestamp 1679581782
transform 1 0 49344 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_515
timestamp 1679581782
transform 1 0 50016 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_522
timestamp 1679581782
transform 1 0 50688 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_529
timestamp 1679581782
transform 1 0 51360 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_536
timestamp 1679581782
transform 1 0 52032 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_543
timestamp 1679581782
transform 1 0 52704 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_550
timestamp 1679581782
transform 1 0 53376 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_557
timestamp 1679581782
transform 1 0 54048 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_564
timestamp 1679581782
transform 1 0 54720 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_571
timestamp 1679581782
transform 1 0 55392 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_578
timestamp 1679581782
transform 1 0 56064 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_585
timestamp 1679581782
transform 1 0 56736 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_592
timestamp 1679581782
transform 1 0 57408 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_599
timestamp 1679581782
transform 1 0 58080 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_606
timestamp 1679581782
transform 1 0 58752 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_613
timestamp 1679581782
transform 1 0 59424 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_620
timestamp 1679581782
transform 1 0 60096 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_627
timestamp 1679581782
transform 1 0 60768 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_634
timestamp 1679581782
transform 1 0 61440 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_641
timestamp 1679581782
transform 1 0 62112 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_648
timestamp 1679581782
transform 1 0 62784 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_655
timestamp 1679581782
transform 1 0 63456 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_662
timestamp 1679581782
transform 1 0 64128 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_669
timestamp 1679581782
transform 1 0 64800 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_676
timestamp 1679581782
transform 1 0 65472 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_683
timestamp 1679581782
transform 1 0 66144 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_690
timestamp 1679581782
transform 1 0 66816 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_697
timestamp 1679581782
transform 1 0 67488 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_704
timestamp 1679581782
transform 1 0 68160 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_711
timestamp 1679581782
transform 1 0 68832 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_718
timestamp 1679581782
transform 1 0 69504 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_725
timestamp 1679581782
transform 1 0 70176 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_732
timestamp 1679581782
transform 1 0 70848 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_739
timestamp 1679581782
transform 1 0 71520 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_746
timestamp 1679581782
transform 1 0 72192 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_753
timestamp 1679581782
transform 1 0 72864 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_760
timestamp 1679581782
transform 1 0 73536 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_767
timestamp 1679581782
transform 1 0 74208 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_774
timestamp 1679581782
transform 1 0 74880 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_781
timestamp 1679581782
transform 1 0 75552 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_788
timestamp 1679581782
transform 1 0 76224 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_795
timestamp 1679581782
transform 1 0 76896 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_802
timestamp 1679581782
transform 1 0 77568 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_809
timestamp 1679581782
transform 1 0 78240 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_816
timestamp 1679581782
transform 1 0 78912 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_823
timestamp 1679581782
transform 1 0 79584 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_830
timestamp 1679581782
transform 1 0 80256 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_837
timestamp 1679581782
transform 1 0 80928 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_844
timestamp 1679581782
transform 1 0 81600 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_851
timestamp 1679581782
transform 1 0 82272 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_858
timestamp 1679581782
transform 1 0 82944 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_865
timestamp 1679581782
transform 1 0 83616 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_872
timestamp 1679581782
transform 1 0 84288 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_879
timestamp 1679581782
transform 1 0 84960 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_886
timestamp 1679581782
transform 1 0 85632 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_893
timestamp 1679581782
transform 1 0 86304 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_900
timestamp 1679581782
transform 1 0 86976 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_907
timestamp 1679581782
transform 1 0 87648 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_914
timestamp 1679581782
transform 1 0 88320 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_921
timestamp 1679581782
transform 1 0 88992 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_928
timestamp 1679581782
transform 1 0 89664 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_935
timestamp 1679581782
transform 1 0 90336 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_942
timestamp 1679581782
transform 1 0 91008 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_949
timestamp 1679581782
transform 1 0 91680 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_956
timestamp 1679581782
transform 1 0 92352 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_963
timestamp 1679581782
transform 1 0 93024 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_970
timestamp 1679581782
transform 1 0 93696 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_977
timestamp 1679581782
transform 1 0 94368 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_984
timestamp 1679581782
transform 1 0 95040 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_991
timestamp 1679581782
transform 1 0 95712 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_998
timestamp 1679581782
transform 1 0 96384 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_1005
timestamp 1679581782
transform 1 0 97056 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_1012
timestamp 1679581782
transform 1 0 97728 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_1019
timestamp 1679581782
transform 1 0 98400 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_1026
timestamp 1677580104
transform 1 0 99072 0 -1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_1028
timestamp 1677579658
transform 1 0 99264 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_4
timestamp 1679581782
transform 1 0 960 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_11
timestamp 1679581782
transform 1 0 1632 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_18
timestamp 1679581782
transform 1 0 2304 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_25
timestamp 1679581782
transform 1 0 2976 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_32
timestamp 1679581782
transform 1 0 3648 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_39
timestamp 1679581782
transform 1 0 4320 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_46
timestamp 1679581782
transform 1 0 4992 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_53
timestamp 1679581782
transform 1 0 5664 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_60
timestamp 1679581782
transform 1 0 6336 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_67
timestamp 1679581782
transform 1 0 7008 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_74
timestamp 1679581782
transform 1 0 7680 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_81
timestamp 1679581782
transform 1 0 8352 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_88
timestamp 1679581782
transform 1 0 9024 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_95
timestamp 1679581782
transform 1 0 9696 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_102
timestamp 1679581782
transform 1 0 10368 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_109
timestamp 1679581782
transform 1 0 11040 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_116
timestamp 1679581782
transform 1 0 11712 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_123
timestamp 1679581782
transform 1 0 12384 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_130
timestamp 1679581782
transform 1 0 13056 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_137
timestamp 1679581782
transform 1 0 13728 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_144
timestamp 1679581782
transform 1 0 14400 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_151
timestamp 1679581782
transform 1 0 15072 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_158
timestamp 1679581782
transform 1 0 15744 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_165
timestamp 1679581782
transform 1 0 16416 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_172
timestamp 1679581782
transform 1 0 17088 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_179
timestamp 1679581782
transform 1 0 17760 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_186
timestamp 1679581782
transform 1 0 18432 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_193
timestamp 1679581782
transform 1 0 19104 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_200
timestamp 1679581782
transform 1 0 19776 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_207
timestamp 1679581782
transform 1 0 20448 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_214
timestamp 1679581782
transform 1 0 21120 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_221
timestamp 1679581782
transform 1 0 21792 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_228
timestamp 1679581782
transform 1 0 22464 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_235
timestamp 1679581782
transform 1 0 23136 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_242
timestamp 1679581782
transform 1 0 23808 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_249
timestamp 1679581782
transform 1 0 24480 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_256
timestamp 1679581782
transform 1 0 25152 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_263
timestamp 1679581782
transform 1 0 25824 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_270
timestamp 1679581782
transform 1 0 26496 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_277
timestamp 1679581782
transform 1 0 27168 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_284
timestamp 1679581782
transform 1 0 27840 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_291
timestamp 1679581782
transform 1 0 28512 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_298
timestamp 1679581782
transform 1 0 29184 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_305
timestamp 1679581782
transform 1 0 29856 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_312
timestamp 1679581782
transform 1 0 30528 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_319
timestamp 1679581782
transform 1 0 31200 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_326
timestamp 1679581782
transform 1 0 31872 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_333
timestamp 1679581782
transform 1 0 32544 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_340
timestamp 1679581782
transform 1 0 33216 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_347
timestamp 1679581782
transform 1 0 33888 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_354
timestamp 1679581782
transform 1 0 34560 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_361
timestamp 1679581782
transform 1 0 35232 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_368
timestamp 1679581782
transform 1 0 35904 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_375
timestamp 1679581782
transform 1 0 36576 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_382
timestamp 1679581782
transform 1 0 37248 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_389
timestamp 1679581782
transform 1 0 37920 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_396
timestamp 1679581782
transform 1 0 38592 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_403
timestamp 1679581782
transform 1 0 39264 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_410
timestamp 1679581782
transform 1 0 39936 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_417
timestamp 1679581782
transform 1 0 40608 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_424
timestamp 1679581782
transform 1 0 41280 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_431
timestamp 1679581782
transform 1 0 41952 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_438
timestamp 1679581782
transform 1 0 42624 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_445
timestamp 1679581782
transform 1 0 43296 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_452
timestamp 1679581782
transform 1 0 43968 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_459
timestamp 1679581782
transform 1 0 44640 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_466
timestamp 1679581782
transform 1 0 45312 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_473
timestamp 1679581782
transform 1 0 45984 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_480
timestamp 1679581782
transform 1 0 46656 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_487
timestamp 1679581782
transform 1 0 47328 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_494
timestamp 1679581782
transform 1 0 48000 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_501
timestamp 1679581782
transform 1 0 48672 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_508
timestamp 1679581782
transform 1 0 49344 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_515
timestamp 1679581782
transform 1 0 50016 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_522
timestamp 1679581782
transform 1 0 50688 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_529
timestamp 1679581782
transform 1 0 51360 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_536
timestamp 1679581782
transform 1 0 52032 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_543
timestamp 1679581782
transform 1 0 52704 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_550
timestamp 1679581782
transform 1 0 53376 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_557
timestamp 1679581782
transform 1 0 54048 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_564
timestamp 1679581782
transform 1 0 54720 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_571
timestamp 1679581782
transform 1 0 55392 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_578
timestamp 1679581782
transform 1 0 56064 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_585
timestamp 1679581782
transform 1 0 56736 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_592
timestamp 1679581782
transform 1 0 57408 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_599
timestamp 1679581782
transform 1 0 58080 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_606
timestamp 1679581782
transform 1 0 58752 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_613
timestamp 1679581782
transform 1 0 59424 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_620
timestamp 1679581782
transform 1 0 60096 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_627
timestamp 1679581782
transform 1 0 60768 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_634
timestamp 1679581782
transform 1 0 61440 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_641
timestamp 1679581782
transform 1 0 62112 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_648
timestamp 1679581782
transform 1 0 62784 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_655
timestamp 1679581782
transform 1 0 63456 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_662
timestamp 1679581782
transform 1 0 64128 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_669
timestamp 1679581782
transform 1 0 64800 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_676
timestamp 1679581782
transform 1 0 65472 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_683
timestamp 1679581782
transform 1 0 66144 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_690
timestamp 1679581782
transform 1 0 66816 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_697
timestamp 1679581782
transform 1 0 67488 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_704
timestamp 1679581782
transform 1 0 68160 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_711
timestamp 1679581782
transform 1 0 68832 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_718
timestamp 1679581782
transform 1 0 69504 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_725
timestamp 1679581782
transform 1 0 70176 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_732
timestamp 1679581782
transform 1 0 70848 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_739
timestamp 1679581782
transform 1 0 71520 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_746
timestamp 1679581782
transform 1 0 72192 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_753
timestamp 1679581782
transform 1 0 72864 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_760
timestamp 1679581782
transform 1 0 73536 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_767
timestamp 1679581782
transform 1 0 74208 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_774
timestamp 1679581782
transform 1 0 74880 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_781
timestamp 1679581782
transform 1 0 75552 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_788
timestamp 1679581782
transform 1 0 76224 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_795
timestamp 1679581782
transform 1 0 76896 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_802
timestamp 1679581782
transform 1 0 77568 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_809
timestamp 1679581782
transform 1 0 78240 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_816
timestamp 1679581782
transform 1 0 78912 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_823
timestamp 1679581782
transform 1 0 79584 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_830
timestamp 1679581782
transform 1 0 80256 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_837
timestamp 1679581782
transform 1 0 80928 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_844
timestamp 1679581782
transform 1 0 81600 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_851
timestamp 1679581782
transform 1 0 82272 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_858
timestamp 1679581782
transform 1 0 82944 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_865
timestamp 1679581782
transform 1 0 83616 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_872
timestamp 1679581782
transform 1 0 84288 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_879
timestamp 1679581782
transform 1 0 84960 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_886
timestamp 1679581782
transform 1 0 85632 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_893
timestamp 1679581782
transform 1 0 86304 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_900
timestamp 1679581782
transform 1 0 86976 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_907
timestamp 1679581782
transform 1 0 87648 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_914
timestamp 1679581782
transform 1 0 88320 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_921
timestamp 1679581782
transform 1 0 88992 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_928
timestamp 1679581782
transform 1 0 89664 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_935
timestamp 1679581782
transform 1 0 90336 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_942
timestamp 1679581782
transform 1 0 91008 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_949
timestamp 1679581782
transform 1 0 91680 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_956
timestamp 1679581782
transform 1 0 92352 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_963
timestamp 1679581782
transform 1 0 93024 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_970
timestamp 1679581782
transform 1 0 93696 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_977
timestamp 1679581782
transform 1 0 94368 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_984
timestamp 1679581782
transform 1 0 95040 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_991
timestamp 1679581782
transform 1 0 95712 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_998
timestamp 1679581782
transform 1 0 96384 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_1005
timestamp 1679581782
transform 1 0 97056 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_1012
timestamp 1679581782
transform 1 0 97728 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_1019
timestamp 1679581782
transform 1 0 98400 0 1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_6_1026
timestamp 1677580104
transform 1 0 99072 0 1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_1028
timestamp 1677579658
transform 1 0 99264 0 1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_0
timestamp 1679581782
transform 1 0 576 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_7
timestamp 1679581782
transform 1 0 1248 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_14
timestamp 1679581782
transform 1 0 1920 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_21
timestamp 1679581782
transform 1 0 2592 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_28
timestamp 1679581782
transform 1 0 3264 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_35
timestamp 1679581782
transform 1 0 3936 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_42
timestamp 1679581782
transform 1 0 4608 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_49
timestamp 1679581782
transform 1 0 5280 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_56
timestamp 1679581782
transform 1 0 5952 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_63
timestamp 1679581782
transform 1 0 6624 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_70
timestamp 1679581782
transform 1 0 7296 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_77
timestamp 1679581782
transform 1 0 7968 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_84
timestamp 1679581782
transform 1 0 8640 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_91
timestamp 1679581782
transform 1 0 9312 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_98
timestamp 1679581782
transform 1 0 9984 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_105
timestamp 1679581782
transform 1 0 10656 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_112
timestamp 1679581782
transform 1 0 11328 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_119
timestamp 1679581782
transform 1 0 12000 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_126
timestamp 1679581782
transform 1 0 12672 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_133
timestamp 1679581782
transform 1 0 13344 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_140
timestamp 1679581782
transform 1 0 14016 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_147
timestamp 1679581782
transform 1 0 14688 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_154
timestamp 1679581782
transform 1 0 15360 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_161
timestamp 1679581782
transform 1 0 16032 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_168
timestamp 1679581782
transform 1 0 16704 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_175
timestamp 1679581782
transform 1 0 17376 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_182
timestamp 1679581782
transform 1 0 18048 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_189
timestamp 1679581782
transform 1 0 18720 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_196
timestamp 1679581782
transform 1 0 19392 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_203
timestamp 1679581782
transform 1 0 20064 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_210
timestamp 1679581782
transform 1 0 20736 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_217
timestamp 1679581782
transform 1 0 21408 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_224
timestamp 1679581782
transform 1 0 22080 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_231
timestamp 1679581782
transform 1 0 22752 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_238
timestamp 1679581782
transform 1 0 23424 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_245
timestamp 1679581782
transform 1 0 24096 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_252
timestamp 1679581782
transform 1 0 24768 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_259
timestamp 1679581782
transform 1 0 25440 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_266
timestamp 1679581782
transform 1 0 26112 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_273
timestamp 1679581782
transform 1 0 26784 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_280
timestamp 1679581782
transform 1 0 27456 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_287
timestamp 1679581782
transform 1 0 28128 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_294
timestamp 1679581782
transform 1 0 28800 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_301
timestamp 1679581782
transform 1 0 29472 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_308
timestamp 1679581782
transform 1 0 30144 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_315
timestamp 1679581782
transform 1 0 30816 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_322
timestamp 1679581782
transform 1 0 31488 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_329
timestamp 1679581782
transform 1 0 32160 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_336
timestamp 1679581782
transform 1 0 32832 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_343
timestamp 1679581782
transform 1 0 33504 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_350
timestamp 1679581782
transform 1 0 34176 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_357
timestamp 1679581782
transform 1 0 34848 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_364
timestamp 1679581782
transform 1 0 35520 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_371
timestamp 1679581782
transform 1 0 36192 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_378
timestamp 1679581782
transform 1 0 36864 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_385
timestamp 1679581782
transform 1 0 37536 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_392
timestamp 1679581782
transform 1 0 38208 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_399
timestamp 1679581782
transform 1 0 38880 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_406
timestamp 1679581782
transform 1 0 39552 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_413
timestamp 1679581782
transform 1 0 40224 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_420
timestamp 1679581782
transform 1 0 40896 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_427
timestamp 1679581782
transform 1 0 41568 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_434
timestamp 1679581782
transform 1 0 42240 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_441
timestamp 1679581782
transform 1 0 42912 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_448
timestamp 1679581782
transform 1 0 43584 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_455
timestamp 1679581782
transform 1 0 44256 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_462
timestamp 1679581782
transform 1 0 44928 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_469
timestamp 1679581782
transform 1 0 45600 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_476
timestamp 1679581782
transform 1 0 46272 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_483
timestamp 1679581782
transform 1 0 46944 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_490
timestamp 1679581782
transform 1 0 47616 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_497
timestamp 1679581782
transform 1 0 48288 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_504
timestamp 1679581782
transform 1 0 48960 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_511
timestamp 1679581782
transform 1 0 49632 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_518
timestamp 1679581782
transform 1 0 50304 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_525
timestamp 1679581782
transform 1 0 50976 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_532
timestamp 1679581782
transform 1 0 51648 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_539
timestamp 1679581782
transform 1 0 52320 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_546
timestamp 1679581782
transform 1 0 52992 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_553
timestamp 1679581782
transform 1 0 53664 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_560
timestamp 1679581782
transform 1 0 54336 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_567
timestamp 1679581782
transform 1 0 55008 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_574
timestamp 1679581782
transform 1 0 55680 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_581
timestamp 1679581782
transform 1 0 56352 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_588
timestamp 1679581782
transform 1 0 57024 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_595
timestamp 1679581782
transform 1 0 57696 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_602
timestamp 1679581782
transform 1 0 58368 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_609
timestamp 1679581782
transform 1 0 59040 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_616
timestamp 1679581782
transform 1 0 59712 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_623
timestamp 1679581782
transform 1 0 60384 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_630
timestamp 1679581782
transform 1 0 61056 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_637
timestamp 1679581782
transform 1 0 61728 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_644
timestamp 1679581782
transform 1 0 62400 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_651
timestamp 1679581782
transform 1 0 63072 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_658
timestamp 1679581782
transform 1 0 63744 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_665
timestamp 1679581782
transform 1 0 64416 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_672
timestamp 1679581782
transform 1 0 65088 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_679
timestamp 1679581782
transform 1 0 65760 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_686
timestamp 1679581782
transform 1 0 66432 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_693
timestamp 1679581782
transform 1 0 67104 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_700
timestamp 1679581782
transform 1 0 67776 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_707
timestamp 1679581782
transform 1 0 68448 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_714
timestamp 1679581782
transform 1 0 69120 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_721
timestamp 1679581782
transform 1 0 69792 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_728
timestamp 1679581782
transform 1 0 70464 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_735
timestamp 1679581782
transform 1 0 71136 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_742
timestamp 1679581782
transform 1 0 71808 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_749
timestamp 1679581782
transform 1 0 72480 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_756
timestamp 1679581782
transform 1 0 73152 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_763
timestamp 1679581782
transform 1 0 73824 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_770
timestamp 1679581782
transform 1 0 74496 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_777
timestamp 1679581782
transform 1 0 75168 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_784
timestamp 1679581782
transform 1 0 75840 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_791
timestamp 1679581782
transform 1 0 76512 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_798
timestamp 1679581782
transform 1 0 77184 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_805
timestamp 1679581782
transform 1 0 77856 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_812
timestamp 1679581782
transform 1 0 78528 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_819
timestamp 1679581782
transform 1 0 79200 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_826
timestamp 1679581782
transform 1 0 79872 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_833
timestamp 1679581782
transform 1 0 80544 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_840
timestamp 1679581782
transform 1 0 81216 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_847
timestamp 1679581782
transform 1 0 81888 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_854
timestamp 1679581782
transform 1 0 82560 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_861
timestamp 1679581782
transform 1 0 83232 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_868
timestamp 1679581782
transform 1 0 83904 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_875
timestamp 1679581782
transform 1 0 84576 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_882
timestamp 1679581782
transform 1 0 85248 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_889
timestamp 1679581782
transform 1 0 85920 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_896
timestamp 1679581782
transform 1 0 86592 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_903
timestamp 1679581782
transform 1 0 87264 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_910
timestamp 1679581782
transform 1 0 87936 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_917
timestamp 1679581782
transform 1 0 88608 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_924
timestamp 1679581782
transform 1 0 89280 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_931
timestamp 1679581782
transform 1 0 89952 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_938
timestamp 1679581782
transform 1 0 90624 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_945
timestamp 1679581782
transform 1 0 91296 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_952
timestamp 1679581782
transform 1 0 91968 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_959
timestamp 1679581782
transform 1 0 92640 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_966
timestamp 1679581782
transform 1 0 93312 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_973
timestamp 1679581782
transform 1 0 93984 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_980
timestamp 1679581782
transform 1 0 94656 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_987
timestamp 1679581782
transform 1 0 95328 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_994
timestamp 1679581782
transform 1 0 96000 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_1001
timestamp 1679581782
transform 1 0 96672 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_1008
timestamp 1679581782
transform 1 0 97344 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_1015
timestamp 1679581782
transform 1 0 98016 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_1022
timestamp 1679581782
transform 1 0 98688 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_4
timestamp 1679581782
transform 1 0 960 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_11
timestamp 1679581782
transform 1 0 1632 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_18
timestamp 1679581782
transform 1 0 2304 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_25
timestamp 1679581782
transform 1 0 2976 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_32
timestamp 1679581782
transform 1 0 3648 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_39
timestamp 1679581782
transform 1 0 4320 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_46
timestamp 1679581782
transform 1 0 4992 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_53
timestamp 1679581782
transform 1 0 5664 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_60
timestamp 1679581782
transform 1 0 6336 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_67
timestamp 1679581782
transform 1 0 7008 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_74
timestamp 1679581782
transform 1 0 7680 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_81
timestamp 1679581782
transform 1 0 8352 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_88
timestamp 1679581782
transform 1 0 9024 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_95
timestamp 1679581782
transform 1 0 9696 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_102
timestamp 1679581782
transform 1 0 10368 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_109
timestamp 1679581782
transform 1 0 11040 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_116
timestamp 1679581782
transform 1 0 11712 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_123
timestamp 1679581782
transform 1 0 12384 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_130
timestamp 1679581782
transform 1 0 13056 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_137
timestamp 1679581782
transform 1 0 13728 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_144
timestamp 1679581782
transform 1 0 14400 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_151
timestamp 1679581782
transform 1 0 15072 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_158
timestamp 1679581782
transform 1 0 15744 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_165
timestamp 1679581782
transform 1 0 16416 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_172
timestamp 1679581782
transform 1 0 17088 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_179
timestamp 1679581782
transform 1 0 17760 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_186
timestamp 1679581782
transform 1 0 18432 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_193
timestamp 1679581782
transform 1 0 19104 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_200
timestamp 1679581782
transform 1 0 19776 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_207
timestamp 1679581782
transform 1 0 20448 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_214
timestamp 1679581782
transform 1 0 21120 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_221
timestamp 1679581782
transform 1 0 21792 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_228
timestamp 1679581782
transform 1 0 22464 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_235
timestamp 1679581782
transform 1 0 23136 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_242
timestamp 1679581782
transform 1 0 23808 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_249
timestamp 1679581782
transform 1 0 24480 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_256
timestamp 1679581782
transform 1 0 25152 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_263
timestamp 1679581782
transform 1 0 25824 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_270
timestamp 1679581782
transform 1 0 26496 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_277
timestamp 1679581782
transform 1 0 27168 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_284
timestamp 1679581782
transform 1 0 27840 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_291
timestamp 1679581782
transform 1 0 28512 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_298
timestamp 1679581782
transform 1 0 29184 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_305
timestamp 1679581782
transform 1 0 29856 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_312
timestamp 1679581782
transform 1 0 30528 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_319
timestamp 1679581782
transform 1 0 31200 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_326
timestamp 1679581782
transform 1 0 31872 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_333
timestamp 1679581782
transform 1 0 32544 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_340
timestamp 1679581782
transform 1 0 33216 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_347
timestamp 1679581782
transform 1 0 33888 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_354
timestamp 1679581782
transform 1 0 34560 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_361
timestamp 1679581782
transform 1 0 35232 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_368
timestamp 1679581782
transform 1 0 35904 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_375
timestamp 1679581782
transform 1 0 36576 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_382
timestamp 1679581782
transform 1 0 37248 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_389
timestamp 1679581782
transform 1 0 37920 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_396
timestamp 1679581782
transform 1 0 38592 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_403
timestamp 1679581782
transform 1 0 39264 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_410
timestamp 1679581782
transform 1 0 39936 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_417
timestamp 1679581782
transform 1 0 40608 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_424
timestamp 1679581782
transform 1 0 41280 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_431
timestamp 1679581782
transform 1 0 41952 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_438
timestamp 1679581782
transform 1 0 42624 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_445
timestamp 1679581782
transform 1 0 43296 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_452
timestamp 1679581782
transform 1 0 43968 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_459
timestamp 1679581782
transform 1 0 44640 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_466
timestamp 1679581782
transform 1 0 45312 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_473
timestamp 1679581782
transform 1 0 45984 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_480
timestamp 1679581782
transform 1 0 46656 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_487
timestamp 1679581782
transform 1 0 47328 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_494
timestamp 1679581782
transform 1 0 48000 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_501
timestamp 1679581782
transform 1 0 48672 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_508
timestamp 1679581782
transform 1 0 49344 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_515
timestamp 1679581782
transform 1 0 50016 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_522
timestamp 1679581782
transform 1 0 50688 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_529
timestamp 1679581782
transform 1 0 51360 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_536
timestamp 1679581782
transform 1 0 52032 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_543
timestamp 1679581782
transform 1 0 52704 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_550
timestamp 1679581782
transform 1 0 53376 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_557
timestamp 1679581782
transform 1 0 54048 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_564
timestamp 1679581782
transform 1 0 54720 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_571
timestamp 1679581782
transform 1 0 55392 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_578
timestamp 1679581782
transform 1 0 56064 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_585
timestamp 1679581782
transform 1 0 56736 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_592
timestamp 1679581782
transform 1 0 57408 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_599
timestamp 1679581782
transform 1 0 58080 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_606
timestamp 1679581782
transform 1 0 58752 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_613
timestamp 1679581782
transform 1 0 59424 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_620
timestamp 1679581782
transform 1 0 60096 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_627
timestamp 1679581782
transform 1 0 60768 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_634
timestamp 1679581782
transform 1 0 61440 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_641
timestamp 1679581782
transform 1 0 62112 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_648
timestamp 1679581782
transform 1 0 62784 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_655
timestamp 1679581782
transform 1 0 63456 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_662
timestamp 1679581782
transform 1 0 64128 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_669
timestamp 1679581782
transform 1 0 64800 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_676
timestamp 1679581782
transform 1 0 65472 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_683
timestamp 1679581782
transform 1 0 66144 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_690
timestamp 1679581782
transform 1 0 66816 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_697
timestamp 1679581782
transform 1 0 67488 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_704
timestamp 1679581782
transform 1 0 68160 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_711
timestamp 1679581782
transform 1 0 68832 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_718
timestamp 1679581782
transform 1 0 69504 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_725
timestamp 1679581782
transform 1 0 70176 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_732
timestamp 1679581782
transform 1 0 70848 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_739
timestamp 1679581782
transform 1 0 71520 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_746
timestamp 1679581782
transform 1 0 72192 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_753
timestamp 1679581782
transform 1 0 72864 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_760
timestamp 1679581782
transform 1 0 73536 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_767
timestamp 1679581782
transform 1 0 74208 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_774
timestamp 1679581782
transform 1 0 74880 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_781
timestamp 1679581782
transform 1 0 75552 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_788
timestamp 1679581782
transform 1 0 76224 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_795
timestamp 1679581782
transform 1 0 76896 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_802
timestamp 1679581782
transform 1 0 77568 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_809
timestamp 1679581782
transform 1 0 78240 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_816
timestamp 1679581782
transform 1 0 78912 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_823
timestamp 1679581782
transform 1 0 79584 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_830
timestamp 1679581782
transform 1 0 80256 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_837
timestamp 1679581782
transform 1 0 80928 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_844
timestamp 1679581782
transform 1 0 81600 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_851
timestamp 1679581782
transform 1 0 82272 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_858
timestamp 1679581782
transform 1 0 82944 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_865
timestamp 1679581782
transform 1 0 83616 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_872
timestamp 1679581782
transform 1 0 84288 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_879
timestamp 1679581782
transform 1 0 84960 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_886
timestamp 1679581782
transform 1 0 85632 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_893
timestamp 1679581782
transform 1 0 86304 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_900
timestamp 1679581782
transform 1 0 86976 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_907
timestamp 1679581782
transform 1 0 87648 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_914
timestamp 1679581782
transform 1 0 88320 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_921
timestamp 1679581782
transform 1 0 88992 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_928
timestamp 1679581782
transform 1 0 89664 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_935
timestamp 1679581782
transform 1 0 90336 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_942
timestamp 1679581782
transform 1 0 91008 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_949
timestamp 1679581782
transform 1 0 91680 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_956
timestamp 1679581782
transform 1 0 92352 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_963
timestamp 1679581782
transform 1 0 93024 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_970
timestamp 1679581782
transform 1 0 93696 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_977
timestamp 1679581782
transform 1 0 94368 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_984
timestamp 1679581782
transform 1 0 95040 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_991
timestamp 1679581782
transform 1 0 95712 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_998
timestamp 1679581782
transform 1 0 96384 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_1005
timestamp 1679581782
transform 1 0 97056 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_1012
timestamp 1679581782
transform 1 0 97728 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_1019
timestamp 1679581782
transform 1 0 98400 0 1 6804
box -48 -56 720 834
use sg13g2_fill_2  FILLER_8_1026
timestamp 1677580104
transform 1 0 99072 0 1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_1028
timestamp 1677579658
transform 1 0 99264 0 1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_4
timestamp 1679581782
transform 1 0 960 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_11
timestamp 1679581782
transform 1 0 1632 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_18
timestamp 1679581782
transform 1 0 2304 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_25
timestamp 1679581782
transform 1 0 2976 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_32
timestamp 1679581782
transform 1 0 3648 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_39
timestamp 1679581782
transform 1 0 4320 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_46
timestamp 1679581782
transform 1 0 4992 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_53
timestamp 1679581782
transform 1 0 5664 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_60
timestamp 1679581782
transform 1 0 6336 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_67
timestamp 1679581782
transform 1 0 7008 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_74
timestamp 1679581782
transform 1 0 7680 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_81
timestamp 1679581782
transform 1 0 8352 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_88
timestamp 1679581782
transform 1 0 9024 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_95
timestamp 1679581782
transform 1 0 9696 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_102
timestamp 1679581782
transform 1 0 10368 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_109
timestamp 1679581782
transform 1 0 11040 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_116
timestamp 1679581782
transform 1 0 11712 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_123
timestamp 1679581782
transform 1 0 12384 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_130
timestamp 1679581782
transform 1 0 13056 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_137
timestamp 1679581782
transform 1 0 13728 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_144
timestamp 1679581782
transform 1 0 14400 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_151
timestamp 1679581782
transform 1 0 15072 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_158
timestamp 1679581782
transform 1 0 15744 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_165
timestamp 1679581782
transform 1 0 16416 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_172
timestamp 1679581782
transform 1 0 17088 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_179
timestamp 1679581782
transform 1 0 17760 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_186
timestamp 1679581782
transform 1 0 18432 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_193
timestamp 1679581782
transform 1 0 19104 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_200
timestamp 1679581782
transform 1 0 19776 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_207
timestamp 1679581782
transform 1 0 20448 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_214
timestamp 1679581782
transform 1 0 21120 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_221
timestamp 1679581782
transform 1 0 21792 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_228
timestamp 1679581782
transform 1 0 22464 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_235
timestamp 1679581782
transform 1 0 23136 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_242
timestamp 1679581782
transform 1 0 23808 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_249
timestamp 1679581782
transform 1 0 24480 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_256
timestamp 1679581782
transform 1 0 25152 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_263
timestamp 1679581782
transform 1 0 25824 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_270
timestamp 1679581782
transform 1 0 26496 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_277
timestamp 1679581782
transform 1 0 27168 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_284
timestamp 1679581782
transform 1 0 27840 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_291
timestamp 1679581782
transform 1 0 28512 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_298
timestamp 1679581782
transform 1 0 29184 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_305
timestamp 1679581782
transform 1 0 29856 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_312
timestamp 1679581782
transform 1 0 30528 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_319
timestamp 1679581782
transform 1 0 31200 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_326
timestamp 1679581782
transform 1 0 31872 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_333
timestamp 1679581782
transform 1 0 32544 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_340
timestamp 1679581782
transform 1 0 33216 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_347
timestamp 1679581782
transform 1 0 33888 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_354
timestamp 1679581782
transform 1 0 34560 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_361
timestamp 1679581782
transform 1 0 35232 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_368
timestamp 1679581782
transform 1 0 35904 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_375
timestamp 1679581782
transform 1 0 36576 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_382
timestamp 1679581782
transform 1 0 37248 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_389
timestamp 1679581782
transform 1 0 37920 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_396
timestamp 1679581782
transform 1 0 38592 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_403
timestamp 1679581782
transform 1 0 39264 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_410
timestamp 1679581782
transform 1 0 39936 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_417
timestamp 1679581782
transform 1 0 40608 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_424
timestamp 1679581782
transform 1 0 41280 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_431
timestamp 1679581782
transform 1 0 41952 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_438
timestamp 1679581782
transform 1 0 42624 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_445
timestamp 1679581782
transform 1 0 43296 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_452
timestamp 1679581782
transform 1 0 43968 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_459
timestamp 1679581782
transform 1 0 44640 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_466
timestamp 1679581782
transform 1 0 45312 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_473
timestamp 1679581782
transform 1 0 45984 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_480
timestamp 1679581782
transform 1 0 46656 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_487
timestamp 1679581782
transform 1 0 47328 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_494
timestamp 1679581782
transform 1 0 48000 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_501
timestamp 1679581782
transform 1 0 48672 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_508
timestamp 1679581782
transform 1 0 49344 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_515
timestamp 1679581782
transform 1 0 50016 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_522
timestamp 1679581782
transform 1 0 50688 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_529
timestamp 1679581782
transform 1 0 51360 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_536
timestamp 1679581782
transform 1 0 52032 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_543
timestamp 1679581782
transform 1 0 52704 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_550
timestamp 1679581782
transform 1 0 53376 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_557
timestamp 1679581782
transform 1 0 54048 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_564
timestamp 1679581782
transform 1 0 54720 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_571
timestamp 1679581782
transform 1 0 55392 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_578
timestamp 1679581782
transform 1 0 56064 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_585
timestamp 1679581782
transform 1 0 56736 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_592
timestamp 1679581782
transform 1 0 57408 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_599
timestamp 1679581782
transform 1 0 58080 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_606
timestamp 1679581782
transform 1 0 58752 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_613
timestamp 1679581782
transform 1 0 59424 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_620
timestamp 1679581782
transform 1 0 60096 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_627
timestamp 1679581782
transform 1 0 60768 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_634
timestamp 1679581782
transform 1 0 61440 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_641
timestamp 1679581782
transform 1 0 62112 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_648
timestamp 1679581782
transform 1 0 62784 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_655
timestamp 1679581782
transform 1 0 63456 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_662
timestamp 1679581782
transform 1 0 64128 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_669
timestamp 1679581782
transform 1 0 64800 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_676
timestamp 1679581782
transform 1 0 65472 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_683
timestamp 1679581782
transform 1 0 66144 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_690
timestamp 1679581782
transform 1 0 66816 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_697
timestamp 1679581782
transform 1 0 67488 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_704
timestamp 1679581782
transform 1 0 68160 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_711
timestamp 1679581782
transform 1 0 68832 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_718
timestamp 1679581782
transform 1 0 69504 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_725
timestamp 1679581782
transform 1 0 70176 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_732
timestamp 1679581782
transform 1 0 70848 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_739
timestamp 1679581782
transform 1 0 71520 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_746
timestamp 1679581782
transform 1 0 72192 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_753
timestamp 1679581782
transform 1 0 72864 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_760
timestamp 1679581782
transform 1 0 73536 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_767
timestamp 1679581782
transform 1 0 74208 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_774
timestamp 1679581782
transform 1 0 74880 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_781
timestamp 1679581782
transform 1 0 75552 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_788
timestamp 1679581782
transform 1 0 76224 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_795
timestamp 1679581782
transform 1 0 76896 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_802
timestamp 1679581782
transform 1 0 77568 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_809
timestamp 1679581782
transform 1 0 78240 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_816
timestamp 1679581782
transform 1 0 78912 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_823
timestamp 1679581782
transform 1 0 79584 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_830
timestamp 1679581782
transform 1 0 80256 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_837
timestamp 1679581782
transform 1 0 80928 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_844
timestamp 1679581782
transform 1 0 81600 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_851
timestamp 1679581782
transform 1 0 82272 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_858
timestamp 1679581782
transform 1 0 82944 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_865
timestamp 1679581782
transform 1 0 83616 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_872
timestamp 1679581782
transform 1 0 84288 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_879
timestamp 1679581782
transform 1 0 84960 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_886
timestamp 1679581782
transform 1 0 85632 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_893
timestamp 1679581782
transform 1 0 86304 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_900
timestamp 1679581782
transform 1 0 86976 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_907
timestamp 1679581782
transform 1 0 87648 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_914
timestamp 1679581782
transform 1 0 88320 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_921
timestamp 1679581782
transform 1 0 88992 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_928
timestamp 1679581782
transform 1 0 89664 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_935
timestamp 1679581782
transform 1 0 90336 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_942
timestamp 1679581782
transform 1 0 91008 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_949
timestamp 1679581782
transform 1 0 91680 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_956
timestamp 1679581782
transform 1 0 92352 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_963
timestamp 1679581782
transform 1 0 93024 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_970
timestamp 1679581782
transform 1 0 93696 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_977
timestamp 1679581782
transform 1 0 94368 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_984
timestamp 1679581782
transform 1 0 95040 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_991
timestamp 1679581782
transform 1 0 95712 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_998
timestamp 1679581782
transform 1 0 96384 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_1005
timestamp 1679581782
transform 1 0 97056 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_1012
timestamp 1679581782
transform 1 0 97728 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_1019
timestamp 1679581782
transform 1 0 98400 0 -1 8316
box -48 -56 720 834
use sg13g2_fill_2  FILLER_9_1026
timestamp 1677580104
transform 1 0 99072 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_1028
timestamp 1677579658
transform 1 0 99264 0 -1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_10_4
timestamp 1679581782
transform 1 0 960 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_11
timestamp 1679581782
transform 1 0 1632 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_18
timestamp 1679581782
transform 1 0 2304 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_25
timestamp 1679581782
transform 1 0 2976 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_32
timestamp 1679581782
transform 1 0 3648 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_39
timestamp 1679581782
transform 1 0 4320 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_46
timestamp 1679581782
transform 1 0 4992 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_53
timestamp 1679581782
transform 1 0 5664 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_60
timestamp 1679581782
transform 1 0 6336 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_67
timestamp 1679581782
transform 1 0 7008 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_74
timestamp 1679581782
transform 1 0 7680 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_81
timestamp 1679581782
transform 1 0 8352 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_88
timestamp 1679581782
transform 1 0 9024 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_95
timestamp 1679581782
transform 1 0 9696 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_102
timestamp 1679581782
transform 1 0 10368 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_109
timestamp 1679581782
transform 1 0 11040 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_116
timestamp 1679581782
transform 1 0 11712 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_123
timestamp 1679581782
transform 1 0 12384 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_130
timestamp 1679581782
transform 1 0 13056 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_137
timestamp 1679581782
transform 1 0 13728 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_144
timestamp 1679581782
transform 1 0 14400 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_151
timestamp 1679581782
transform 1 0 15072 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_158
timestamp 1679581782
transform 1 0 15744 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_165
timestamp 1679581782
transform 1 0 16416 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_172
timestamp 1679581782
transform 1 0 17088 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_179
timestamp 1679581782
transform 1 0 17760 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_186
timestamp 1679581782
transform 1 0 18432 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_193
timestamp 1679581782
transform 1 0 19104 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_200
timestamp 1679581782
transform 1 0 19776 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_207
timestamp 1679581782
transform 1 0 20448 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_214
timestamp 1679581782
transform 1 0 21120 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_221
timestamp 1679581782
transform 1 0 21792 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_228
timestamp 1679581782
transform 1 0 22464 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_235
timestamp 1679581782
transform 1 0 23136 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_242
timestamp 1679581782
transform 1 0 23808 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_249
timestamp 1679581782
transform 1 0 24480 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_256
timestamp 1679581782
transform 1 0 25152 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_263
timestamp 1679581782
transform 1 0 25824 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_270
timestamp 1679581782
transform 1 0 26496 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_277
timestamp 1679581782
transform 1 0 27168 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_284
timestamp 1679581782
transform 1 0 27840 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_291
timestamp 1679581782
transform 1 0 28512 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_298
timestamp 1679581782
transform 1 0 29184 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_305
timestamp 1679581782
transform 1 0 29856 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_312
timestamp 1679581782
transform 1 0 30528 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_319
timestamp 1679581782
transform 1 0 31200 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_326
timestamp 1679581782
transform 1 0 31872 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_333
timestamp 1679581782
transform 1 0 32544 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_340
timestamp 1679581782
transform 1 0 33216 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_347
timestamp 1679581782
transform 1 0 33888 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_354
timestamp 1679581782
transform 1 0 34560 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_361
timestamp 1679581782
transform 1 0 35232 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_368
timestamp 1679581782
transform 1 0 35904 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_375
timestamp 1679581782
transform 1 0 36576 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_382
timestamp 1679581782
transform 1 0 37248 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_389
timestamp 1679581782
transform 1 0 37920 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_396
timestamp 1679581782
transform 1 0 38592 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_403
timestamp 1679581782
transform 1 0 39264 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_410
timestamp 1679581782
transform 1 0 39936 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_417
timestamp 1679581782
transform 1 0 40608 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_424
timestamp 1679581782
transform 1 0 41280 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_431
timestamp 1679581782
transform 1 0 41952 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_438
timestamp 1679581782
transform 1 0 42624 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_445
timestamp 1679581782
transform 1 0 43296 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_452
timestamp 1679581782
transform 1 0 43968 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_459
timestamp 1679581782
transform 1 0 44640 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_466
timestamp 1679581782
transform 1 0 45312 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_473
timestamp 1679581782
transform 1 0 45984 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_480
timestamp 1679581782
transform 1 0 46656 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_487
timestamp 1679581782
transform 1 0 47328 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_494
timestamp 1679581782
transform 1 0 48000 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_501
timestamp 1679581782
transform 1 0 48672 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_508
timestamp 1679581782
transform 1 0 49344 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_515
timestamp 1679581782
transform 1 0 50016 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_522
timestamp 1679581782
transform 1 0 50688 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_529
timestamp 1679581782
transform 1 0 51360 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_536
timestamp 1679581782
transform 1 0 52032 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_543
timestamp 1679581782
transform 1 0 52704 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_550
timestamp 1679581782
transform 1 0 53376 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_557
timestamp 1679581782
transform 1 0 54048 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_564
timestamp 1679581782
transform 1 0 54720 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_571
timestamp 1679581782
transform 1 0 55392 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_578
timestamp 1679581782
transform 1 0 56064 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_585
timestamp 1679581782
transform 1 0 56736 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_592
timestamp 1679581782
transform 1 0 57408 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_599
timestamp 1679581782
transform 1 0 58080 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_606
timestamp 1679581782
transform 1 0 58752 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_613
timestamp 1679581782
transform 1 0 59424 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_620
timestamp 1679581782
transform 1 0 60096 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_627
timestamp 1679581782
transform 1 0 60768 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_634
timestamp 1679581782
transform 1 0 61440 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_641
timestamp 1679581782
transform 1 0 62112 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_648
timestamp 1679581782
transform 1 0 62784 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_655
timestamp 1679581782
transform 1 0 63456 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_662
timestamp 1679581782
transform 1 0 64128 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_669
timestamp 1679581782
transform 1 0 64800 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_676
timestamp 1679581782
transform 1 0 65472 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_683
timestamp 1679581782
transform 1 0 66144 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_690
timestamp 1679581782
transform 1 0 66816 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_697
timestamp 1679581782
transform 1 0 67488 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_704
timestamp 1679581782
transform 1 0 68160 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_711
timestamp 1679581782
transform 1 0 68832 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_718
timestamp 1679581782
transform 1 0 69504 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_725
timestamp 1679581782
transform 1 0 70176 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_732
timestamp 1679581782
transform 1 0 70848 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_739
timestamp 1679581782
transform 1 0 71520 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_746
timestamp 1679581782
transform 1 0 72192 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_753
timestamp 1679581782
transform 1 0 72864 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_760
timestamp 1679581782
transform 1 0 73536 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_767
timestamp 1679581782
transform 1 0 74208 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_774
timestamp 1679581782
transform 1 0 74880 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_781
timestamp 1679581782
transform 1 0 75552 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_788
timestamp 1679581782
transform 1 0 76224 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_795
timestamp 1679581782
transform 1 0 76896 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_802
timestamp 1679581782
transform 1 0 77568 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_809
timestamp 1679581782
transform 1 0 78240 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_816
timestamp 1679581782
transform 1 0 78912 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_823
timestamp 1679581782
transform 1 0 79584 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_830
timestamp 1679581782
transform 1 0 80256 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_837
timestamp 1679581782
transform 1 0 80928 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_844
timestamp 1679581782
transform 1 0 81600 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_851
timestamp 1679581782
transform 1 0 82272 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_858
timestamp 1679581782
transform 1 0 82944 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_865
timestamp 1679581782
transform 1 0 83616 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_872
timestamp 1679581782
transform 1 0 84288 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_879
timestamp 1679581782
transform 1 0 84960 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_886
timestamp 1679581782
transform 1 0 85632 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_893
timestamp 1679581782
transform 1 0 86304 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_900
timestamp 1679581782
transform 1 0 86976 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_907
timestamp 1679581782
transform 1 0 87648 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_914
timestamp 1679581782
transform 1 0 88320 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_921
timestamp 1679581782
transform 1 0 88992 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_928
timestamp 1679581782
transform 1 0 89664 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_935
timestamp 1679581782
transform 1 0 90336 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_942
timestamp 1679581782
transform 1 0 91008 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_949
timestamp 1679581782
transform 1 0 91680 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_956
timestamp 1679581782
transform 1 0 92352 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_963
timestamp 1679581782
transform 1 0 93024 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_970
timestamp 1679581782
transform 1 0 93696 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_977
timestamp 1679581782
transform 1 0 94368 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_984
timestamp 1679581782
transform 1 0 95040 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_991
timestamp 1679581782
transform 1 0 95712 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_998
timestamp 1679581782
transform 1 0 96384 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_1005
timestamp 1679581782
transform 1 0 97056 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_1012
timestamp 1679581782
transform 1 0 97728 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_1019
timestamp 1679581782
transform 1 0 98400 0 1 8316
box -48 -56 720 834
use sg13g2_fill_2  FILLER_10_1026
timestamp 1677580104
transform 1 0 99072 0 1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_1028
timestamp 1677579658
transform 1 0 99264 0 1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_11_4
timestamp 1679581782
transform 1 0 960 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_11
timestamp 1679581782
transform 1 0 1632 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_18
timestamp 1679581782
transform 1 0 2304 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_25
timestamp 1679581782
transform 1 0 2976 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_32
timestamp 1679581782
transform 1 0 3648 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_39
timestamp 1679581782
transform 1 0 4320 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_46
timestamp 1679581782
transform 1 0 4992 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_53
timestamp 1679581782
transform 1 0 5664 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_60
timestamp 1679581782
transform 1 0 6336 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_67
timestamp 1679581782
transform 1 0 7008 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_74
timestamp 1679581782
transform 1 0 7680 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_81
timestamp 1679581782
transform 1 0 8352 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_88
timestamp 1679581782
transform 1 0 9024 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_95
timestamp 1679581782
transform 1 0 9696 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_102
timestamp 1679581782
transform 1 0 10368 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_109
timestamp 1679581782
transform 1 0 11040 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_116
timestamp 1679581782
transform 1 0 11712 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_123
timestamp 1679581782
transform 1 0 12384 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_130
timestamp 1679581782
transform 1 0 13056 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_137
timestamp 1679581782
transform 1 0 13728 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_144
timestamp 1679581782
transform 1 0 14400 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_151
timestamp 1679581782
transform 1 0 15072 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_158
timestamp 1679581782
transform 1 0 15744 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_165
timestamp 1679581782
transform 1 0 16416 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_172
timestamp 1679581782
transform 1 0 17088 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_179
timestamp 1679581782
transform 1 0 17760 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_186
timestamp 1679581782
transform 1 0 18432 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_193
timestamp 1679581782
transform 1 0 19104 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_200
timestamp 1679581782
transform 1 0 19776 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_207
timestamp 1679581782
transform 1 0 20448 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_214
timestamp 1679581782
transform 1 0 21120 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_221
timestamp 1679581782
transform 1 0 21792 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_228
timestamp 1679581782
transform 1 0 22464 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_235
timestamp 1679581782
transform 1 0 23136 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_242
timestamp 1679581782
transform 1 0 23808 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_249
timestamp 1679581782
transform 1 0 24480 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_256
timestamp 1679581782
transform 1 0 25152 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_263
timestamp 1679581782
transform 1 0 25824 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_270
timestamp 1679581782
transform 1 0 26496 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_277
timestamp 1679581782
transform 1 0 27168 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_284
timestamp 1679581782
transform 1 0 27840 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_291
timestamp 1679581782
transform 1 0 28512 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_298
timestamp 1679581782
transform 1 0 29184 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_305
timestamp 1679581782
transform 1 0 29856 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_312
timestamp 1679581782
transform 1 0 30528 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_319
timestamp 1679581782
transform 1 0 31200 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_326
timestamp 1679581782
transform 1 0 31872 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_333
timestamp 1679581782
transform 1 0 32544 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_340
timestamp 1679581782
transform 1 0 33216 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_347
timestamp 1679581782
transform 1 0 33888 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_354
timestamp 1679581782
transform 1 0 34560 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_361
timestamp 1679581782
transform 1 0 35232 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_368
timestamp 1679581782
transform 1 0 35904 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_375
timestamp 1679581782
transform 1 0 36576 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_382
timestamp 1679581782
transform 1 0 37248 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_389
timestamp 1679581782
transform 1 0 37920 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_396
timestamp 1679581782
transform 1 0 38592 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_403
timestamp 1679581782
transform 1 0 39264 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_410
timestamp 1679581782
transform 1 0 39936 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_417
timestamp 1679581782
transform 1 0 40608 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_424
timestamp 1679581782
transform 1 0 41280 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_431
timestamp 1679581782
transform 1 0 41952 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_438
timestamp 1679581782
transform 1 0 42624 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_445
timestamp 1679581782
transform 1 0 43296 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_452
timestamp 1679581782
transform 1 0 43968 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_459
timestamp 1679581782
transform 1 0 44640 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_466
timestamp 1679581782
transform 1 0 45312 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_473
timestamp 1679581782
transform 1 0 45984 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_480
timestamp 1679581782
transform 1 0 46656 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_487
timestamp 1679581782
transform 1 0 47328 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_494
timestamp 1679581782
transform 1 0 48000 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_501
timestamp 1679581782
transform 1 0 48672 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_508
timestamp 1679581782
transform 1 0 49344 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_515
timestamp 1679581782
transform 1 0 50016 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_522
timestamp 1679581782
transform 1 0 50688 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_529
timestamp 1679581782
transform 1 0 51360 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_536
timestamp 1679581782
transform 1 0 52032 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_543
timestamp 1679581782
transform 1 0 52704 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_550
timestamp 1679581782
transform 1 0 53376 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_557
timestamp 1679581782
transform 1 0 54048 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_564
timestamp 1679581782
transform 1 0 54720 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_571
timestamp 1679581782
transform 1 0 55392 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_578
timestamp 1679581782
transform 1 0 56064 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_585
timestamp 1679581782
transform 1 0 56736 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_592
timestamp 1679581782
transform 1 0 57408 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_599
timestamp 1679581782
transform 1 0 58080 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_606
timestamp 1679581782
transform 1 0 58752 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_613
timestamp 1679581782
transform 1 0 59424 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_620
timestamp 1679581782
transform 1 0 60096 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_627
timestamp 1679581782
transform 1 0 60768 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_634
timestamp 1679581782
transform 1 0 61440 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_641
timestamp 1679581782
transform 1 0 62112 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_648
timestamp 1679581782
transform 1 0 62784 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_655
timestamp 1679581782
transform 1 0 63456 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_662
timestamp 1679581782
transform 1 0 64128 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_669
timestamp 1679581782
transform 1 0 64800 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_676
timestamp 1679581782
transform 1 0 65472 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_683
timestamp 1679581782
transform 1 0 66144 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_690
timestamp 1679581782
transform 1 0 66816 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_697
timestamp 1679581782
transform 1 0 67488 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_704
timestamp 1679581782
transform 1 0 68160 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_711
timestamp 1679581782
transform 1 0 68832 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_718
timestamp 1679581782
transform 1 0 69504 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_725
timestamp 1679581782
transform 1 0 70176 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_732
timestamp 1679581782
transform 1 0 70848 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_739
timestamp 1679581782
transform 1 0 71520 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_746
timestamp 1679581782
transform 1 0 72192 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_753
timestamp 1679581782
transform 1 0 72864 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_760
timestamp 1679581782
transform 1 0 73536 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_767
timestamp 1679581782
transform 1 0 74208 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_774
timestamp 1679581782
transform 1 0 74880 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_781
timestamp 1679581782
transform 1 0 75552 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_788
timestamp 1679581782
transform 1 0 76224 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_795
timestamp 1679581782
transform 1 0 76896 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_802
timestamp 1679581782
transform 1 0 77568 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_809
timestamp 1679581782
transform 1 0 78240 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_816
timestamp 1679581782
transform 1 0 78912 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_823
timestamp 1679581782
transform 1 0 79584 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_830
timestamp 1679581782
transform 1 0 80256 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_837
timestamp 1679581782
transform 1 0 80928 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_844
timestamp 1679581782
transform 1 0 81600 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_851
timestamp 1679581782
transform 1 0 82272 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_858
timestamp 1679581782
transform 1 0 82944 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_865
timestamp 1679581782
transform 1 0 83616 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_872
timestamp 1679581782
transform 1 0 84288 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_879
timestamp 1679581782
transform 1 0 84960 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_886
timestamp 1679581782
transform 1 0 85632 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_893
timestamp 1679581782
transform 1 0 86304 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_900
timestamp 1679581782
transform 1 0 86976 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_907
timestamp 1679581782
transform 1 0 87648 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_914
timestamp 1679581782
transform 1 0 88320 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_921
timestamp 1679581782
transform 1 0 88992 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_928
timestamp 1679581782
transform 1 0 89664 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_935
timestamp 1679581782
transform 1 0 90336 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_942
timestamp 1679581782
transform 1 0 91008 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_949
timestamp 1679581782
transform 1 0 91680 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_956
timestamp 1679581782
transform 1 0 92352 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_963
timestamp 1679581782
transform 1 0 93024 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_970
timestamp 1679581782
transform 1 0 93696 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_977
timestamp 1679581782
transform 1 0 94368 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_984
timestamp 1679581782
transform 1 0 95040 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_991
timestamp 1679581782
transform 1 0 95712 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_998
timestamp 1679581782
transform 1 0 96384 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_1005
timestamp 1679581782
transform 1 0 97056 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_1012
timestamp 1679581782
transform 1 0 97728 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_1019
timestamp 1679581782
transform 1 0 98400 0 -1 9828
box -48 -56 720 834
use sg13g2_fill_2  FILLER_11_1026
timestamp 1677580104
transform 1 0 99072 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_1028
timestamp 1677579658
transform 1 0 99264 0 -1 9828
box -48 -56 144 834
use sg13g2_decap_8  FILLER_12_4
timestamp 1679581782
transform 1 0 960 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_11
timestamp 1679581782
transform 1 0 1632 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_18
timestamp 1679581782
transform 1 0 2304 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_25
timestamp 1679581782
transform 1 0 2976 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_32
timestamp 1679581782
transform 1 0 3648 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_39
timestamp 1679581782
transform 1 0 4320 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_46
timestamp 1679581782
transform 1 0 4992 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_53
timestamp 1679581782
transform 1 0 5664 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_60
timestamp 1679581782
transform 1 0 6336 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_67
timestamp 1679581782
transform 1 0 7008 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_74
timestamp 1679581782
transform 1 0 7680 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_81
timestamp 1679581782
transform 1 0 8352 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_88
timestamp 1679581782
transform 1 0 9024 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_95
timestamp 1679581782
transform 1 0 9696 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_102
timestamp 1679581782
transform 1 0 10368 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_109
timestamp 1679581782
transform 1 0 11040 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_116
timestamp 1679581782
transform 1 0 11712 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_123
timestamp 1679581782
transform 1 0 12384 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_130
timestamp 1679581782
transform 1 0 13056 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_137
timestamp 1679581782
transform 1 0 13728 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_144
timestamp 1679581782
transform 1 0 14400 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_151
timestamp 1679581782
transform 1 0 15072 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_158
timestamp 1679581782
transform 1 0 15744 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_165
timestamp 1679581782
transform 1 0 16416 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_172
timestamp 1679581782
transform 1 0 17088 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_179
timestamp 1679581782
transform 1 0 17760 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_186
timestamp 1679581782
transform 1 0 18432 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_193
timestamp 1679581782
transform 1 0 19104 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_200
timestamp 1679581782
transform 1 0 19776 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_207
timestamp 1679581782
transform 1 0 20448 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_214
timestamp 1679581782
transform 1 0 21120 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_221
timestamp 1679581782
transform 1 0 21792 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_228
timestamp 1679581782
transform 1 0 22464 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_235
timestamp 1679581782
transform 1 0 23136 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_242
timestamp 1679581782
transform 1 0 23808 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_249
timestamp 1679581782
transform 1 0 24480 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_256
timestamp 1679581782
transform 1 0 25152 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_263
timestamp 1679581782
transform 1 0 25824 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_270
timestamp 1679581782
transform 1 0 26496 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_277
timestamp 1679581782
transform 1 0 27168 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_284
timestamp 1679581782
transform 1 0 27840 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_291
timestamp 1679581782
transform 1 0 28512 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_298
timestamp 1679581782
transform 1 0 29184 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_305
timestamp 1679581782
transform 1 0 29856 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_312
timestamp 1679581782
transform 1 0 30528 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_319
timestamp 1679581782
transform 1 0 31200 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_326
timestamp 1679581782
transform 1 0 31872 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_333
timestamp 1679581782
transform 1 0 32544 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_340
timestamp 1679581782
transform 1 0 33216 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_347
timestamp 1679581782
transform 1 0 33888 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_354
timestamp 1679581782
transform 1 0 34560 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_361
timestamp 1679581782
transform 1 0 35232 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_368
timestamp 1679581782
transform 1 0 35904 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_375
timestamp 1679581782
transform 1 0 36576 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_382
timestamp 1679581782
transform 1 0 37248 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_389
timestamp 1679581782
transform 1 0 37920 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_396
timestamp 1679581782
transform 1 0 38592 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_403
timestamp 1679581782
transform 1 0 39264 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_410
timestamp 1679581782
transform 1 0 39936 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_417
timestamp 1679581782
transform 1 0 40608 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_424
timestamp 1679581782
transform 1 0 41280 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_431
timestamp 1679581782
transform 1 0 41952 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_438
timestamp 1679581782
transform 1 0 42624 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_445
timestamp 1679581782
transform 1 0 43296 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_452
timestamp 1679581782
transform 1 0 43968 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_459
timestamp 1679581782
transform 1 0 44640 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_466
timestamp 1679581782
transform 1 0 45312 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_473
timestamp 1679581782
transform 1 0 45984 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_480
timestamp 1679581782
transform 1 0 46656 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_487
timestamp 1679581782
transform 1 0 47328 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_494
timestamp 1679581782
transform 1 0 48000 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_501
timestamp 1679581782
transform 1 0 48672 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_508
timestamp 1679581782
transform 1 0 49344 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_515
timestamp 1679581782
transform 1 0 50016 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_522
timestamp 1679581782
transform 1 0 50688 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_529
timestamp 1679581782
transform 1 0 51360 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_536
timestamp 1679581782
transform 1 0 52032 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_543
timestamp 1679581782
transform 1 0 52704 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_550
timestamp 1679581782
transform 1 0 53376 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_557
timestamp 1679581782
transform 1 0 54048 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_564
timestamp 1679581782
transform 1 0 54720 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_571
timestamp 1679581782
transform 1 0 55392 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_578
timestamp 1679581782
transform 1 0 56064 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_585
timestamp 1679581782
transform 1 0 56736 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_592
timestamp 1679581782
transform 1 0 57408 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_599
timestamp 1679581782
transform 1 0 58080 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_606
timestamp 1679581782
transform 1 0 58752 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_613
timestamp 1679581782
transform 1 0 59424 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_620
timestamp 1679581782
transform 1 0 60096 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_627
timestamp 1679581782
transform 1 0 60768 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_634
timestamp 1679581782
transform 1 0 61440 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_641
timestamp 1679581782
transform 1 0 62112 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_648
timestamp 1679581782
transform 1 0 62784 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_655
timestamp 1679581782
transform 1 0 63456 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_662
timestamp 1679581782
transform 1 0 64128 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_669
timestamp 1679581782
transform 1 0 64800 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_676
timestamp 1679581782
transform 1 0 65472 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_683
timestamp 1679581782
transform 1 0 66144 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_690
timestamp 1679581782
transform 1 0 66816 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_697
timestamp 1679581782
transform 1 0 67488 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_704
timestamp 1679581782
transform 1 0 68160 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_711
timestamp 1679581782
transform 1 0 68832 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_718
timestamp 1679581782
transform 1 0 69504 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_725
timestamp 1679581782
transform 1 0 70176 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_732
timestamp 1679581782
transform 1 0 70848 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_739
timestamp 1679581782
transform 1 0 71520 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_746
timestamp 1679581782
transform 1 0 72192 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_753
timestamp 1679581782
transform 1 0 72864 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_760
timestamp 1679581782
transform 1 0 73536 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_767
timestamp 1679581782
transform 1 0 74208 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_774
timestamp 1679581782
transform 1 0 74880 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_781
timestamp 1679581782
transform 1 0 75552 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_788
timestamp 1679581782
transform 1 0 76224 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_795
timestamp 1679581782
transform 1 0 76896 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_802
timestamp 1679581782
transform 1 0 77568 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_809
timestamp 1679581782
transform 1 0 78240 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_816
timestamp 1679581782
transform 1 0 78912 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_823
timestamp 1679581782
transform 1 0 79584 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_830
timestamp 1679581782
transform 1 0 80256 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_837
timestamp 1679581782
transform 1 0 80928 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_844
timestamp 1679581782
transform 1 0 81600 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_851
timestamp 1679581782
transform 1 0 82272 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_858
timestamp 1679581782
transform 1 0 82944 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_865
timestamp 1679581782
transform 1 0 83616 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_872
timestamp 1679581782
transform 1 0 84288 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_879
timestamp 1679581782
transform 1 0 84960 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_886
timestamp 1679581782
transform 1 0 85632 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_893
timestamp 1679581782
transform 1 0 86304 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_900
timestamp 1679581782
transform 1 0 86976 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_907
timestamp 1679581782
transform 1 0 87648 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_914
timestamp 1679581782
transform 1 0 88320 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_921
timestamp 1679581782
transform 1 0 88992 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_928
timestamp 1679581782
transform 1 0 89664 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_935
timestamp 1679581782
transform 1 0 90336 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_942
timestamp 1679581782
transform 1 0 91008 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_949
timestamp 1679581782
transform 1 0 91680 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_956
timestamp 1679581782
transform 1 0 92352 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_963
timestamp 1679581782
transform 1 0 93024 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_970
timestamp 1679581782
transform 1 0 93696 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_977
timestamp 1679581782
transform 1 0 94368 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_984
timestamp 1679581782
transform 1 0 95040 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_991
timestamp 1679581782
transform 1 0 95712 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_998
timestamp 1679581782
transform 1 0 96384 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_1005
timestamp 1679581782
transform 1 0 97056 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_1012
timestamp 1679581782
transform 1 0 97728 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_1019
timestamp 1679581782
transform 1 0 98400 0 1 9828
box -48 -56 720 834
use sg13g2_fill_2  FILLER_12_1026
timestamp 1677580104
transform 1 0 99072 0 1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_12_1028
timestamp 1677579658
transform 1 0 99264 0 1 9828
box -48 -56 144 834
use sg13g2_decap_8  FILLER_13_4
timestamp 1679581782
transform 1 0 960 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_11
timestamp 1679581782
transform 1 0 1632 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_18
timestamp 1679581782
transform 1 0 2304 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_25
timestamp 1679581782
transform 1 0 2976 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_32
timestamp 1679581782
transform 1 0 3648 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_39
timestamp 1679581782
transform 1 0 4320 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_46
timestamp 1679581782
transform 1 0 4992 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_53
timestamp 1679581782
transform 1 0 5664 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_60
timestamp 1679581782
transform 1 0 6336 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_67
timestamp 1679581782
transform 1 0 7008 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_74
timestamp 1679581782
transform 1 0 7680 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_81
timestamp 1679581782
transform 1 0 8352 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_88
timestamp 1679581782
transform 1 0 9024 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_95
timestamp 1679581782
transform 1 0 9696 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_102
timestamp 1679581782
transform 1 0 10368 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_109
timestamp 1679581782
transform 1 0 11040 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_116
timestamp 1679581782
transform 1 0 11712 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_123
timestamp 1679581782
transform 1 0 12384 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_130
timestamp 1679581782
transform 1 0 13056 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_137
timestamp 1679581782
transform 1 0 13728 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_144
timestamp 1679581782
transform 1 0 14400 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_151
timestamp 1679581782
transform 1 0 15072 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_158
timestamp 1679581782
transform 1 0 15744 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_165
timestamp 1679581782
transform 1 0 16416 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_172
timestamp 1679581782
transform 1 0 17088 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_179
timestamp 1679581782
transform 1 0 17760 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_186
timestamp 1679581782
transform 1 0 18432 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_193
timestamp 1679581782
transform 1 0 19104 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_200
timestamp 1679581782
transform 1 0 19776 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_207
timestamp 1679581782
transform 1 0 20448 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_214
timestamp 1679581782
transform 1 0 21120 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_221
timestamp 1679581782
transform 1 0 21792 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_228
timestamp 1679581782
transform 1 0 22464 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_235
timestamp 1679581782
transform 1 0 23136 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_242
timestamp 1679581782
transform 1 0 23808 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_249
timestamp 1679581782
transform 1 0 24480 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_256
timestamp 1679581782
transform 1 0 25152 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_263
timestamp 1679581782
transform 1 0 25824 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_270
timestamp 1679581782
transform 1 0 26496 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_277
timestamp 1679581782
transform 1 0 27168 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_284
timestamp 1679581782
transform 1 0 27840 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_291
timestamp 1679581782
transform 1 0 28512 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_298
timestamp 1679581782
transform 1 0 29184 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_305
timestamp 1679581782
transform 1 0 29856 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_312
timestamp 1679581782
transform 1 0 30528 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_319
timestamp 1679581782
transform 1 0 31200 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_326
timestamp 1679581782
transform 1 0 31872 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_333
timestamp 1679581782
transform 1 0 32544 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_340
timestamp 1679581782
transform 1 0 33216 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_347
timestamp 1679581782
transform 1 0 33888 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_354
timestamp 1679581782
transform 1 0 34560 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_361
timestamp 1679581782
transform 1 0 35232 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_368
timestamp 1679581782
transform 1 0 35904 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_375
timestamp 1679581782
transform 1 0 36576 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_382
timestamp 1679581782
transform 1 0 37248 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_389
timestamp 1679581782
transform 1 0 37920 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_396
timestamp 1679581782
transform 1 0 38592 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_403
timestamp 1679581782
transform 1 0 39264 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_410
timestamp 1679581782
transform 1 0 39936 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_417
timestamp 1679581782
transform 1 0 40608 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_424
timestamp 1679581782
transform 1 0 41280 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_431
timestamp 1679581782
transform 1 0 41952 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_438
timestamp 1679581782
transform 1 0 42624 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_445
timestamp 1679581782
transform 1 0 43296 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_452
timestamp 1679581782
transform 1 0 43968 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_459
timestamp 1679581782
transform 1 0 44640 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_466
timestamp 1679581782
transform 1 0 45312 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_473
timestamp 1679581782
transform 1 0 45984 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_480
timestamp 1679581782
transform 1 0 46656 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_487
timestamp 1679581782
transform 1 0 47328 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_494
timestamp 1679581782
transform 1 0 48000 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_501
timestamp 1679581782
transform 1 0 48672 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_508
timestamp 1679581782
transform 1 0 49344 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_515
timestamp 1679581782
transform 1 0 50016 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_522
timestamp 1679581782
transform 1 0 50688 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_529
timestamp 1679581782
transform 1 0 51360 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_536
timestamp 1679581782
transform 1 0 52032 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_543
timestamp 1679581782
transform 1 0 52704 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_550
timestamp 1679581782
transform 1 0 53376 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_557
timestamp 1679581782
transform 1 0 54048 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_564
timestamp 1679581782
transform 1 0 54720 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_571
timestamp 1679581782
transform 1 0 55392 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_578
timestamp 1679581782
transform 1 0 56064 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_585
timestamp 1679581782
transform 1 0 56736 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_592
timestamp 1679581782
transform 1 0 57408 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_599
timestamp 1679581782
transform 1 0 58080 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_606
timestamp 1679581782
transform 1 0 58752 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_613
timestamp 1679581782
transform 1 0 59424 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_620
timestamp 1679581782
transform 1 0 60096 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_627
timestamp 1679581782
transform 1 0 60768 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_634
timestamp 1679581782
transform 1 0 61440 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_641
timestamp 1679581782
transform 1 0 62112 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_648
timestamp 1679581782
transform 1 0 62784 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_655
timestamp 1679581782
transform 1 0 63456 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_662
timestamp 1679581782
transform 1 0 64128 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_669
timestamp 1679581782
transform 1 0 64800 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_676
timestamp 1679581782
transform 1 0 65472 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_683
timestamp 1679581782
transform 1 0 66144 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_690
timestamp 1679581782
transform 1 0 66816 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_697
timestamp 1679581782
transform 1 0 67488 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_704
timestamp 1679581782
transform 1 0 68160 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_711
timestamp 1679581782
transform 1 0 68832 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_718
timestamp 1679581782
transform 1 0 69504 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_725
timestamp 1679581782
transform 1 0 70176 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_732
timestamp 1679581782
transform 1 0 70848 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_739
timestamp 1679581782
transform 1 0 71520 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_746
timestamp 1679581782
transform 1 0 72192 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_753
timestamp 1679581782
transform 1 0 72864 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_760
timestamp 1679581782
transform 1 0 73536 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_767
timestamp 1679581782
transform 1 0 74208 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_774
timestamp 1679581782
transform 1 0 74880 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_781
timestamp 1679581782
transform 1 0 75552 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_788
timestamp 1679581782
transform 1 0 76224 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_795
timestamp 1679581782
transform 1 0 76896 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_802
timestamp 1679581782
transform 1 0 77568 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_809
timestamp 1679581782
transform 1 0 78240 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_816
timestamp 1679581782
transform 1 0 78912 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_823
timestamp 1679581782
transform 1 0 79584 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_830
timestamp 1679581782
transform 1 0 80256 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_837
timestamp 1679581782
transform 1 0 80928 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_844
timestamp 1679581782
transform 1 0 81600 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_851
timestamp 1679581782
transform 1 0 82272 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_858
timestamp 1679581782
transform 1 0 82944 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_865
timestamp 1679581782
transform 1 0 83616 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_872
timestamp 1679581782
transform 1 0 84288 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_879
timestamp 1679581782
transform 1 0 84960 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_886
timestamp 1679581782
transform 1 0 85632 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_893
timestamp 1679581782
transform 1 0 86304 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_900
timestamp 1679581782
transform 1 0 86976 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_907
timestamp 1679581782
transform 1 0 87648 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_914
timestamp 1679581782
transform 1 0 88320 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_921
timestamp 1679581782
transform 1 0 88992 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_928
timestamp 1679581782
transform 1 0 89664 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_935
timestamp 1679581782
transform 1 0 90336 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_942
timestamp 1679581782
transform 1 0 91008 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_949
timestamp 1679581782
transform 1 0 91680 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_956
timestamp 1679581782
transform 1 0 92352 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_963
timestamp 1679581782
transform 1 0 93024 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_970
timestamp 1679581782
transform 1 0 93696 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_977
timestamp 1679581782
transform 1 0 94368 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_984
timestamp 1679581782
transform 1 0 95040 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_991
timestamp 1679581782
transform 1 0 95712 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_998
timestamp 1679581782
transform 1 0 96384 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_1005
timestamp 1679581782
transform 1 0 97056 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_1012
timestamp 1679581782
transform 1 0 97728 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_1019
timestamp 1679581782
transform 1 0 98400 0 -1 11340
box -48 -56 720 834
use sg13g2_fill_2  FILLER_13_1026
timestamp 1677580104
transform 1 0 99072 0 -1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_13_1028
timestamp 1677579658
transform 1 0 99264 0 -1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_14_4
timestamp 1679581782
transform 1 0 960 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_11
timestamp 1679581782
transform 1 0 1632 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_18
timestamp 1679581782
transform 1 0 2304 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_25
timestamp 1679581782
transform 1 0 2976 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_32
timestamp 1679581782
transform 1 0 3648 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_39
timestamp 1679581782
transform 1 0 4320 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_46
timestamp 1679581782
transform 1 0 4992 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_53
timestamp 1679581782
transform 1 0 5664 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_60
timestamp 1679581782
transform 1 0 6336 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_67
timestamp 1679581782
transform 1 0 7008 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_74
timestamp 1679581782
transform 1 0 7680 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_81
timestamp 1679581782
transform 1 0 8352 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_88
timestamp 1679581782
transform 1 0 9024 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_95
timestamp 1679581782
transform 1 0 9696 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_102
timestamp 1679581782
transform 1 0 10368 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_109
timestamp 1679581782
transform 1 0 11040 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_116
timestamp 1679581782
transform 1 0 11712 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_123
timestamp 1679581782
transform 1 0 12384 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_130
timestamp 1679581782
transform 1 0 13056 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_137
timestamp 1679581782
transform 1 0 13728 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_144
timestamp 1679581782
transform 1 0 14400 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_151
timestamp 1679581782
transform 1 0 15072 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_158
timestamp 1679581782
transform 1 0 15744 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_165
timestamp 1679581782
transform 1 0 16416 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_172
timestamp 1679581782
transform 1 0 17088 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_179
timestamp 1679581782
transform 1 0 17760 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_186
timestamp 1679581782
transform 1 0 18432 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_193
timestamp 1679581782
transform 1 0 19104 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_200
timestamp 1679581782
transform 1 0 19776 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_207
timestamp 1679581782
transform 1 0 20448 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_214
timestamp 1679581782
transform 1 0 21120 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_221
timestamp 1679581782
transform 1 0 21792 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_255
timestamp 1679581782
transform 1 0 25056 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_262
timestamp 1679581782
transform 1 0 25728 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_269
timestamp 1679581782
transform 1 0 26400 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_276
timestamp 1679581782
transform 1 0 27072 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_283
timestamp 1679581782
transform 1 0 27744 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_290
timestamp 1679581782
transform 1 0 28416 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_297
timestamp 1679581782
transform 1 0 29088 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_304
timestamp 1679581782
transform 1 0 29760 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_311
timestamp 1679581782
transform 1 0 30432 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_318
timestamp 1679581782
transform 1 0 31104 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_325
timestamp 1679581782
transform 1 0 31776 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_332
timestamp 1679581782
transform 1 0 32448 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_339
timestamp 1679581782
transform 1 0 33120 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_346
timestamp 1679581782
transform 1 0 33792 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_353
timestamp 1679581782
transform 1 0 34464 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_360
timestamp 1679581782
transform 1 0 35136 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_367
timestamp 1679581782
transform 1 0 35808 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_374
timestamp 1679581782
transform 1 0 36480 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_381
timestamp 1679581782
transform 1 0 37152 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_388
timestamp 1679581782
transform 1 0 37824 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_395
timestamp 1679581782
transform 1 0 38496 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_402
timestamp 1679581782
transform 1 0 39168 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_409
timestamp 1679581782
transform 1 0 39840 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_416
timestamp 1679581782
transform 1 0 40512 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_423
timestamp 1679581782
transform 1 0 41184 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_430
timestamp 1679581782
transform 1 0 41856 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_437
timestamp 1679581782
transform 1 0 42528 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_444
timestamp 1679581782
transform 1 0 43200 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_451
timestamp 1679581782
transform 1 0 43872 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_458
timestamp 1679581782
transform 1 0 44544 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_465
timestamp 1679581782
transform 1 0 45216 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_472
timestamp 1679581782
transform 1 0 45888 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_479
timestamp 1679581782
transform 1 0 46560 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_486
timestamp 1679581782
transform 1 0 47232 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_493
timestamp 1679581782
transform 1 0 47904 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_500
timestamp 1679581782
transform 1 0 48576 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_507
timestamp 1679581782
transform 1 0 49248 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_514
timestamp 1679581782
transform 1 0 49920 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_521
timestamp 1679581782
transform 1 0 50592 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_528
timestamp 1679581782
transform 1 0 51264 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_535
timestamp 1679581782
transform 1 0 51936 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_542
timestamp 1679581782
transform 1 0 52608 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_549
timestamp 1679581782
transform 1 0 53280 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_556
timestamp 1679581782
transform 1 0 53952 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_563
timestamp 1679581782
transform 1 0 54624 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_570
timestamp 1679581782
transform 1 0 55296 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_577
timestamp 1679581782
transform 1 0 55968 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_584
timestamp 1679581782
transform 1 0 56640 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_591
timestamp 1679581782
transform 1 0 57312 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_598
timestamp 1679581782
transform 1 0 57984 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_605
timestamp 1679581782
transform 1 0 58656 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_612
timestamp 1679581782
transform 1 0 59328 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_619
timestamp 1679581782
transform 1 0 60000 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_626
timestamp 1679581782
transform 1 0 60672 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_633
timestamp 1679581782
transform 1 0 61344 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_640
timestamp 1679581782
transform 1 0 62016 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_647
timestamp 1679581782
transform 1 0 62688 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_654
timestamp 1679581782
transform 1 0 63360 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_661
timestamp 1679581782
transform 1 0 64032 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_668
timestamp 1679581782
transform 1 0 64704 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_675
timestamp 1679581782
transform 1 0 65376 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_682
timestamp 1679581782
transform 1 0 66048 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_689
timestamp 1679581782
transform 1 0 66720 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_696
timestamp 1679581782
transform 1 0 67392 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_703
timestamp 1679581782
transform 1 0 68064 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_710
timestamp 1679581782
transform 1 0 68736 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_717
timestamp 1679581782
transform 1 0 69408 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_724
timestamp 1679581782
transform 1 0 70080 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_731
timestamp 1679581782
transform 1 0 70752 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_738
timestamp 1679581782
transform 1 0 71424 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_745
timestamp 1679581782
transform 1 0 72096 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_752
timestamp 1679581782
transform 1 0 72768 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_759
timestamp 1679581782
transform 1 0 73440 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_766
timestamp 1679581782
transform 1 0 74112 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_773
timestamp 1679581782
transform 1 0 74784 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_780
timestamp 1679581782
transform 1 0 75456 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_787
timestamp 1679581782
transform 1 0 76128 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_794
timestamp 1679581782
transform 1 0 76800 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_801
timestamp 1679581782
transform 1 0 77472 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_808
timestamp 1679581782
transform 1 0 78144 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_815
timestamp 1679581782
transform 1 0 78816 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_822
timestamp 1679581782
transform 1 0 79488 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_829
timestamp 1679581782
transform 1 0 80160 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_836
timestamp 1679581782
transform 1 0 80832 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_843
timestamp 1679581782
transform 1 0 81504 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_850
timestamp 1679581782
transform 1 0 82176 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_857
timestamp 1679581782
transform 1 0 82848 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_864
timestamp 1679581782
transform 1 0 83520 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_871
timestamp 1679581782
transform 1 0 84192 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_878
timestamp 1679581782
transform 1 0 84864 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_885
timestamp 1679581782
transform 1 0 85536 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_892
timestamp 1679581782
transform 1 0 86208 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_899
timestamp 1679581782
transform 1 0 86880 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_906
timestamp 1679581782
transform 1 0 87552 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_913
timestamp 1679581782
transform 1 0 88224 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_920
timestamp 1679581782
transform 1 0 88896 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_927
timestamp 1679581782
transform 1 0 89568 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_934
timestamp 1679581782
transform 1 0 90240 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_941
timestamp 1679581782
transform 1 0 90912 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_948
timestamp 1679581782
transform 1 0 91584 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_955
timestamp 1679581782
transform 1 0 92256 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_962
timestamp 1679581782
transform 1 0 92928 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_969
timestamp 1679581782
transform 1 0 93600 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_976
timestamp 1679581782
transform 1 0 94272 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_983
timestamp 1679581782
transform 1 0 94944 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_990
timestamp 1679581782
transform 1 0 95616 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_997
timestamp 1679581782
transform 1 0 96288 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_1004
timestamp 1679581782
transform 1 0 96960 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_1011
timestamp 1679581782
transform 1 0 97632 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_1018
timestamp 1679581782
transform 1 0 98304 0 1 11340
box -48 -56 720 834
use sg13g2_decap_4  FILLER_14_1025
timestamp 1679577901
transform 1 0 98976 0 1 11340
box -48 -56 432 834
use sg13g2_decap_8  FILLER_15_4
timestamp 1679581782
transform 1 0 960 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_11
timestamp 1679581782
transform 1 0 1632 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_18
timestamp 1679581782
transform 1 0 2304 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_25
timestamp 1679581782
transform 1 0 2976 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_32
timestamp 1679581782
transform 1 0 3648 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_39
timestamp 1679581782
transform 1 0 4320 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_46
timestamp 1679581782
transform 1 0 4992 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_53
timestamp 1679581782
transform 1 0 5664 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_60
timestamp 1679581782
transform 1 0 6336 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_67
timestamp 1679581782
transform 1 0 7008 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_74
timestamp 1679581782
transform 1 0 7680 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_81
timestamp 1679581782
transform 1 0 8352 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_88
timestamp 1679581782
transform 1 0 9024 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_95
timestamp 1679581782
transform 1 0 9696 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_102
timestamp 1679581782
transform 1 0 10368 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_109
timestamp 1679581782
transform 1 0 11040 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_116
timestamp 1679581782
transform 1 0 11712 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_123
timestamp 1679581782
transform 1 0 12384 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_130
timestamp 1679581782
transform 1 0 13056 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_137
timestamp 1679581782
transform 1 0 13728 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_144
timestamp 1679581782
transform 1 0 14400 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_151
timestamp 1679581782
transform 1 0 15072 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_158
timestamp 1679581782
transform 1 0 15744 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_165
timestamp 1679581782
transform 1 0 16416 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_4  FILLER_15_172
timestamp 1679577901
transform 1 0 17088 0 -1 12852
box -48 -56 432 834
use sg13g2_fill_2  FILLER_15_176
timestamp 1677580104
transform 1 0 17472 0 -1 12852
box -48 -56 240 834
use sg13g2_decap_8  FILLER_15_205
timestamp 1679581782
transform 1 0 20256 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_212
timestamp 1679581782
transform 1 0 20928 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_219
timestamp 1679581782
transform 1 0 21600 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_226
timestamp 1679581782
transform 1 0 22272 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_233
timestamp 1679581782
transform 1 0 22944 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_240
timestamp 1679581782
transform 1 0 23616 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_247
timestamp 1679581782
transform 1 0 24288 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_254
timestamp 1679581782
transform 1 0 24960 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_261
timestamp 1679581782
transform 1 0 25632 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_288
timestamp 1679581782
transform 1 0 28224 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_295
timestamp 1679581782
transform 1 0 28896 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_302
timestamp 1679581782
transform 1 0 29568 0 -1 12852
box -48 -56 720 834
use sg13g2_fill_2  FILLER_15_309
timestamp 1677580104
transform 1 0 30240 0 -1 12852
box -48 -56 240 834
use sg13g2_decap_8  FILLER_15_343
timestamp 1679581782
transform 1 0 33504 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_350
timestamp 1679581782
transform 1 0 34176 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_357
timestamp 1679581782
transform 1 0 34848 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_364
timestamp 1679581782
transform 1 0 35520 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_371
timestamp 1679581782
transform 1 0 36192 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_378
timestamp 1679581782
transform 1 0 36864 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_385
timestamp 1679581782
transform 1 0 37536 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_392
timestamp 1679581782
transform 1 0 38208 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_399
timestamp 1679581782
transform 1 0 38880 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_406
timestamp 1679581782
transform 1 0 39552 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_413
timestamp 1679581782
transform 1 0 40224 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_420
timestamp 1679581782
transform 1 0 40896 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_427
timestamp 1679581782
transform 1 0 41568 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_434
timestamp 1679581782
transform 1 0 42240 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_441
timestamp 1679581782
transform 1 0 42912 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_448
timestamp 1679581782
transform 1 0 43584 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_455
timestamp 1679581782
transform 1 0 44256 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_462
timestamp 1679581782
transform 1 0 44928 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_469
timestamp 1679581782
transform 1 0 45600 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_476
timestamp 1679581782
transform 1 0 46272 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_483
timestamp 1679581782
transform 1 0 46944 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_490
timestamp 1679581782
transform 1 0 47616 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_497
timestamp 1679581782
transform 1 0 48288 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_504
timestamp 1679581782
transform 1 0 48960 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_511
timestamp 1679581782
transform 1 0 49632 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_518
timestamp 1679581782
transform 1 0 50304 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_525
timestamp 1679581782
transform 1 0 50976 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_532
timestamp 1679581782
transform 1 0 51648 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_539
timestamp 1679581782
transform 1 0 52320 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_546
timestamp 1679581782
transform 1 0 52992 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_553
timestamp 1679581782
transform 1 0 53664 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_560
timestamp 1679581782
transform 1 0 54336 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_567
timestamp 1679581782
transform 1 0 55008 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_574
timestamp 1679581782
transform 1 0 55680 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_581
timestamp 1679581782
transform 1 0 56352 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_588
timestamp 1679581782
transform 1 0 57024 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_595
timestamp 1679581782
transform 1 0 57696 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_602
timestamp 1679581782
transform 1 0 58368 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_609
timestamp 1679581782
transform 1 0 59040 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_616
timestamp 1679581782
transform 1 0 59712 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_623
timestamp 1679581782
transform 1 0 60384 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_630
timestamp 1679581782
transform 1 0 61056 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_637
timestamp 1679581782
transform 1 0 61728 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_644
timestamp 1679581782
transform 1 0 62400 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_651
timestamp 1679581782
transform 1 0 63072 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_658
timestamp 1679581782
transform 1 0 63744 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_665
timestamp 1679581782
transform 1 0 64416 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_672
timestamp 1679581782
transform 1 0 65088 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_679
timestamp 1679581782
transform 1 0 65760 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_686
timestamp 1679581782
transform 1 0 66432 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_693
timestamp 1679581782
transform 1 0 67104 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_700
timestamp 1679581782
transform 1 0 67776 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_707
timestamp 1679581782
transform 1 0 68448 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_714
timestamp 1679581782
transform 1 0 69120 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_721
timestamp 1679581782
transform 1 0 69792 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_728
timestamp 1679581782
transform 1 0 70464 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_735
timestamp 1679581782
transform 1 0 71136 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_742
timestamp 1679581782
transform 1 0 71808 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_749
timestamp 1679581782
transform 1 0 72480 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_756
timestamp 1679581782
transform 1 0 73152 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_763
timestamp 1679581782
transform 1 0 73824 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_770
timestamp 1679581782
transform 1 0 74496 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_777
timestamp 1679581782
transform 1 0 75168 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_784
timestamp 1679581782
transform 1 0 75840 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_791
timestamp 1679581782
transform 1 0 76512 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_798
timestamp 1679581782
transform 1 0 77184 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_805
timestamp 1679581782
transform 1 0 77856 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_812
timestamp 1679581782
transform 1 0 78528 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_819
timestamp 1679581782
transform 1 0 79200 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_826
timestamp 1679581782
transform 1 0 79872 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_833
timestamp 1679581782
transform 1 0 80544 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_840
timestamp 1679581782
transform 1 0 81216 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_847
timestamp 1679581782
transform 1 0 81888 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_854
timestamp 1679581782
transform 1 0 82560 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_861
timestamp 1679581782
transform 1 0 83232 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_868
timestamp 1679581782
transform 1 0 83904 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_875
timestamp 1679581782
transform 1 0 84576 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_882
timestamp 1679581782
transform 1 0 85248 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_889
timestamp 1679581782
transform 1 0 85920 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_896
timestamp 1679581782
transform 1 0 86592 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_903
timestamp 1679581782
transform 1 0 87264 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_910
timestamp 1679581782
transform 1 0 87936 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_917
timestamp 1679581782
transform 1 0 88608 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_924
timestamp 1679581782
transform 1 0 89280 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_931
timestamp 1679581782
transform 1 0 89952 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_938
timestamp 1679581782
transform 1 0 90624 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_945
timestamp 1679581782
transform 1 0 91296 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_952
timestamp 1679581782
transform 1 0 91968 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_959
timestamp 1679581782
transform 1 0 92640 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_966
timestamp 1679581782
transform 1 0 93312 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_973
timestamp 1679581782
transform 1 0 93984 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_980
timestamp 1679581782
transform 1 0 94656 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_987
timestamp 1679581782
transform 1 0 95328 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_994
timestamp 1679581782
transform 1 0 96000 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_1001
timestamp 1679581782
transform 1 0 96672 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_1008
timestamp 1679581782
transform 1 0 97344 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_1015
timestamp 1679581782
transform 1 0 98016 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_1022
timestamp 1679581782
transform 1 0 98688 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_4
timestamp 1679581782
transform 1 0 960 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_11
timestamp 1679581782
transform 1 0 1632 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_18
timestamp 1679581782
transform 1 0 2304 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_25
timestamp 1679581782
transform 1 0 2976 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_32
timestamp 1679581782
transform 1 0 3648 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_39
timestamp 1679581782
transform 1 0 4320 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_46
timestamp 1679581782
transform 1 0 4992 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_53
timestamp 1679581782
transform 1 0 5664 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_60
timestamp 1679581782
transform 1 0 6336 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_67
timestamp 1679581782
transform 1 0 7008 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_74
timestamp 1679581782
transform 1 0 7680 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_81
timestamp 1679581782
transform 1 0 8352 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_88
timestamp 1679581782
transform 1 0 9024 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_95
timestamp 1679581782
transform 1 0 9696 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_102
timestamp 1679581782
transform 1 0 10368 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_109
timestamp 1679581782
transform 1 0 11040 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_116
timestamp 1679581782
transform 1 0 11712 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_123
timestamp 1679581782
transform 1 0 12384 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_130
timestamp 1679581782
transform 1 0 13056 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_137
timestamp 1679581782
transform 1 0 13728 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_144
timestamp 1679581782
transform 1 0 14400 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_151
timestamp 1679581782
transform 1 0 15072 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_158
timestamp 1679581782
transform 1 0 15744 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_165
timestamp 1679581782
transform 1 0 16416 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_172
timestamp 1679581782
transform 1 0 17088 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_179
timestamp 1679581782
transform 1 0 17760 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_186
timestamp 1679581782
transform 1 0 18432 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_193
timestamp 1679581782
transform 1 0 19104 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_200
timestamp 1679581782
transform 1 0 19776 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_207
timestamp 1679581782
transform 1 0 20448 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_214
timestamp 1679581782
transform 1 0 21120 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_221
timestamp 1679581782
transform 1 0 21792 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_228
timestamp 1679581782
transform 1 0 22464 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_235
timestamp 1679581782
transform 1 0 23136 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_242
timestamp 1679581782
transform 1 0 23808 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_249
timestamp 1679581782
transform 1 0 24480 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_256
timestamp 1679581782
transform 1 0 25152 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_263
timestamp 1679581782
transform 1 0 25824 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_270
timestamp 1679581782
transform 1 0 26496 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_277
timestamp 1679581782
transform 1 0 27168 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_284
timestamp 1679581782
transform 1 0 27840 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_291
timestamp 1679581782
transform 1 0 28512 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_298
timestamp 1679581782
transform 1 0 29184 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_305
timestamp 1679581782
transform 1 0 29856 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_312
timestamp 1679581782
transform 1 0 30528 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_319
timestamp 1679581782
transform 1 0 31200 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_326
timestamp 1679581782
transform 1 0 31872 0 1 12852
box -48 -56 720 834
use sg13g2_decap_4  FILLER_16_333
timestamp 1679577901
transform 1 0 32544 0 1 12852
box -48 -56 432 834
use sg13g2_decap_8  FILLER_16_342
timestamp 1679581782
transform 1 0 33408 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_349
timestamp 1679581782
transform 1 0 34080 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_356
timestamp 1679581782
transform 1 0 34752 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_363
timestamp 1679581782
transform 1 0 35424 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_370
timestamp 1679581782
transform 1 0 36096 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_377
timestamp 1679581782
transform 1 0 36768 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_384
timestamp 1679581782
transform 1 0 37440 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_391
timestamp 1679581782
transform 1 0 38112 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_398
timestamp 1679581782
transform 1 0 38784 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_405
timestamp 1679581782
transform 1 0 39456 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_412
timestamp 1679581782
transform 1 0 40128 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_419
timestamp 1679581782
transform 1 0 40800 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_426
timestamp 1679581782
transform 1 0 41472 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_433
timestamp 1679581782
transform 1 0 42144 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_440
timestamp 1679581782
transform 1 0 42816 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_447
timestamp 1679581782
transform 1 0 43488 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_454
timestamp 1679581782
transform 1 0 44160 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_461
timestamp 1679581782
transform 1 0 44832 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_468
timestamp 1679581782
transform 1 0 45504 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_475
timestamp 1679581782
transform 1 0 46176 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_482
timestamp 1679581782
transform 1 0 46848 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_489
timestamp 1679581782
transform 1 0 47520 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_496
timestamp 1679581782
transform 1 0 48192 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_503
timestamp 1679581782
transform 1 0 48864 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_510
timestamp 1679581782
transform 1 0 49536 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_517
timestamp 1679581782
transform 1 0 50208 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_524
timestamp 1679581782
transform 1 0 50880 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_531
timestamp 1679581782
transform 1 0 51552 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_538
timestamp 1679581782
transform 1 0 52224 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_545
timestamp 1679581782
transform 1 0 52896 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_552
timestamp 1679581782
transform 1 0 53568 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_559
timestamp 1679581782
transform 1 0 54240 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_566
timestamp 1679581782
transform 1 0 54912 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_573
timestamp 1679581782
transform 1 0 55584 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_580
timestamp 1679581782
transform 1 0 56256 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_587
timestamp 1679581782
transform 1 0 56928 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_594
timestamp 1679581782
transform 1 0 57600 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_601
timestamp 1679581782
transform 1 0 58272 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_608
timestamp 1679581782
transform 1 0 58944 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_615
timestamp 1679581782
transform 1 0 59616 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_622
timestamp 1679581782
transform 1 0 60288 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_629
timestamp 1679581782
transform 1 0 60960 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_636
timestamp 1679581782
transform 1 0 61632 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_643
timestamp 1679581782
transform 1 0 62304 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_650
timestamp 1679581782
transform 1 0 62976 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_657
timestamp 1679581782
transform 1 0 63648 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_664
timestamp 1679581782
transform 1 0 64320 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_671
timestamp 1679581782
transform 1 0 64992 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_678
timestamp 1679581782
transform 1 0 65664 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_685
timestamp 1679581782
transform 1 0 66336 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_692
timestamp 1679581782
transform 1 0 67008 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_699
timestamp 1679581782
transform 1 0 67680 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_706
timestamp 1679581782
transform 1 0 68352 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_713
timestamp 1679581782
transform 1 0 69024 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_720
timestamp 1679581782
transform 1 0 69696 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_727
timestamp 1679581782
transform 1 0 70368 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_734
timestamp 1679581782
transform 1 0 71040 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_741
timestamp 1679581782
transform 1 0 71712 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_748
timestamp 1679581782
transform 1 0 72384 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_755
timestamp 1679581782
transform 1 0 73056 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_762
timestamp 1679581782
transform 1 0 73728 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_769
timestamp 1679581782
transform 1 0 74400 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_776
timestamp 1679581782
transform 1 0 75072 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_783
timestamp 1679581782
transform 1 0 75744 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_790
timestamp 1679581782
transform 1 0 76416 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_797
timestamp 1679581782
transform 1 0 77088 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_804
timestamp 1679581782
transform 1 0 77760 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_811
timestamp 1679581782
transform 1 0 78432 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_818
timestamp 1679581782
transform 1 0 79104 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_825
timestamp 1679581782
transform 1 0 79776 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_832
timestamp 1679581782
transform 1 0 80448 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_839
timestamp 1679581782
transform 1 0 81120 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_846
timestamp 1679581782
transform 1 0 81792 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_853
timestamp 1679581782
transform 1 0 82464 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_860
timestamp 1679581782
transform 1 0 83136 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_867
timestamp 1679581782
transform 1 0 83808 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_874
timestamp 1679581782
transform 1 0 84480 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_881
timestamp 1679581782
transform 1 0 85152 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_888
timestamp 1679581782
transform 1 0 85824 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_895
timestamp 1679581782
transform 1 0 86496 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_902
timestamp 1679581782
transform 1 0 87168 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_909
timestamp 1679581782
transform 1 0 87840 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_916
timestamp 1679581782
transform 1 0 88512 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_923
timestamp 1679581782
transform 1 0 89184 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_930
timestamp 1679581782
transform 1 0 89856 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_937
timestamp 1679581782
transform 1 0 90528 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_944
timestamp 1679581782
transform 1 0 91200 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_951
timestamp 1679581782
transform 1 0 91872 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_958
timestamp 1679581782
transform 1 0 92544 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_965
timestamp 1679581782
transform 1 0 93216 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_972
timestamp 1679581782
transform 1 0 93888 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_979
timestamp 1679581782
transform 1 0 94560 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_986
timestamp 1679581782
transform 1 0 95232 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_993
timestamp 1679581782
transform 1 0 95904 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_1000
timestamp 1679581782
transform 1 0 96576 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_1007
timestamp 1679581782
transform 1 0 97248 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_1014
timestamp 1679581782
transform 1 0 97920 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_1021
timestamp 1679581782
transform 1 0 98592 0 1 12852
box -48 -56 720 834
use sg13g2_fill_1  FILLER_16_1028
timestamp 1677579658
transform 1 0 99264 0 1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_17_0
timestamp 1679581782
transform 1 0 576 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_7
timestamp 1679581782
transform 1 0 1248 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_14
timestamp 1679581782
transform 1 0 1920 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_21
timestamp 1679581782
transform 1 0 2592 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_28
timestamp 1679581782
transform 1 0 3264 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_35
timestamp 1679581782
transform 1 0 3936 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_42
timestamp 1679581782
transform 1 0 4608 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_49
timestamp 1679581782
transform 1 0 5280 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_56
timestamp 1679581782
transform 1 0 5952 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_63
timestamp 1679581782
transform 1 0 6624 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_70
timestamp 1679581782
transform 1 0 7296 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_77
timestamp 1679581782
transform 1 0 7968 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_84
timestamp 1679581782
transform 1 0 8640 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_91
timestamp 1679581782
transform 1 0 9312 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_98
timestamp 1679581782
transform 1 0 9984 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_105
timestamp 1679581782
transform 1 0 10656 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_112
timestamp 1679581782
transform 1 0 11328 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_119
timestamp 1679581782
transform 1 0 12000 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_126
timestamp 1679581782
transform 1 0 12672 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_133
timestamp 1679581782
transform 1 0 13344 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_140
timestamp 1679581782
transform 1 0 14016 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_147
timestamp 1679581782
transform 1 0 14688 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_154
timestamp 1679581782
transform 1 0 15360 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_161
timestamp 1679581782
transform 1 0 16032 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_168
timestamp 1679581782
transform 1 0 16704 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_175
timestamp 1679581782
transform 1 0 17376 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_182
timestamp 1679581782
transform 1 0 18048 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_189
timestamp 1679581782
transform 1 0 18720 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_196
timestamp 1679581782
transform 1 0 19392 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_203
timestamp 1679581782
transform 1 0 20064 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_210
timestamp 1679581782
transform 1 0 20736 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_217
timestamp 1679581782
transform 1 0 21408 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_224
timestamp 1679581782
transform 1 0 22080 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_231
timestamp 1679581782
transform 1 0 22752 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_238
timestamp 1679581782
transform 1 0 23424 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_245
timestamp 1679581782
transform 1 0 24096 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_252
timestamp 1679581782
transform 1 0 24768 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_259
timestamp 1679581782
transform 1 0 25440 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_266
timestamp 1679581782
transform 1 0 26112 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_273
timestamp 1679581782
transform 1 0 26784 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_280
timestamp 1679581782
transform 1 0 27456 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_287
timestamp 1679581782
transform 1 0 28128 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_294
timestamp 1679581782
transform 1 0 28800 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_301
timestamp 1679581782
transform 1 0 29472 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_308
timestamp 1679581782
transform 1 0 30144 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_315
timestamp 1679581782
transform 1 0 30816 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_322
timestamp 1679581782
transform 1 0 31488 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_329
timestamp 1679581782
transform 1 0 32160 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_336
timestamp 1679581782
transform 1 0 32832 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_343
timestamp 1679581782
transform 1 0 33504 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_350
timestamp 1679581782
transform 1 0 34176 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_357
timestamp 1679581782
transform 1 0 34848 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_364
timestamp 1679581782
transform 1 0 35520 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_371
timestamp 1679581782
transform 1 0 36192 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_378
timestamp 1679581782
transform 1 0 36864 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_385
timestamp 1679581782
transform 1 0 37536 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_392
timestamp 1679581782
transform 1 0 38208 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_399
timestamp 1679581782
transform 1 0 38880 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_406
timestamp 1679581782
transform 1 0 39552 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_413
timestamp 1679581782
transform 1 0 40224 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_420
timestamp 1679581782
transform 1 0 40896 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_427
timestamp 1679581782
transform 1 0 41568 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_434
timestamp 1679581782
transform 1 0 42240 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_441
timestamp 1679581782
transform 1 0 42912 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_448
timestamp 1679581782
transform 1 0 43584 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_455
timestamp 1679581782
transform 1 0 44256 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_462
timestamp 1679581782
transform 1 0 44928 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_469
timestamp 1679581782
transform 1 0 45600 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_476
timestamp 1679581782
transform 1 0 46272 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_483
timestamp 1679581782
transform 1 0 46944 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_490
timestamp 1679581782
transform 1 0 47616 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_497
timestamp 1679581782
transform 1 0 48288 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_504
timestamp 1679581782
transform 1 0 48960 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_511
timestamp 1679581782
transform 1 0 49632 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_518
timestamp 1679581782
transform 1 0 50304 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_525
timestamp 1679581782
transform 1 0 50976 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_532
timestamp 1679581782
transform 1 0 51648 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_539
timestamp 1679581782
transform 1 0 52320 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_546
timestamp 1679581782
transform 1 0 52992 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_553
timestamp 1679581782
transform 1 0 53664 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_560
timestamp 1679581782
transform 1 0 54336 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_567
timestamp 1679581782
transform 1 0 55008 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_574
timestamp 1679581782
transform 1 0 55680 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_581
timestamp 1679581782
transform 1 0 56352 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_588
timestamp 1679581782
transform 1 0 57024 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_595
timestamp 1679581782
transform 1 0 57696 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_602
timestamp 1679581782
transform 1 0 58368 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_609
timestamp 1679581782
transform 1 0 59040 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_616
timestamp 1679581782
transform 1 0 59712 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_623
timestamp 1679581782
transform 1 0 60384 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_630
timestamp 1679581782
transform 1 0 61056 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_637
timestamp 1679581782
transform 1 0 61728 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_644
timestamp 1679581782
transform 1 0 62400 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_651
timestamp 1679581782
transform 1 0 63072 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_658
timestamp 1679581782
transform 1 0 63744 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_665
timestamp 1679581782
transform 1 0 64416 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_672
timestamp 1679581782
transform 1 0 65088 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_679
timestamp 1679581782
transform 1 0 65760 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_686
timestamp 1679581782
transform 1 0 66432 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_693
timestamp 1679581782
transform 1 0 67104 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_700
timestamp 1679581782
transform 1 0 67776 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_707
timestamp 1679581782
transform 1 0 68448 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_714
timestamp 1679581782
transform 1 0 69120 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_721
timestamp 1679581782
transform 1 0 69792 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_728
timestamp 1679581782
transform 1 0 70464 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_735
timestamp 1679581782
transform 1 0 71136 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_742
timestamp 1679581782
transform 1 0 71808 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_749
timestamp 1679581782
transform 1 0 72480 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_756
timestamp 1679581782
transform 1 0 73152 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_763
timestamp 1679581782
transform 1 0 73824 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_770
timestamp 1679581782
transform 1 0 74496 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_777
timestamp 1679581782
transform 1 0 75168 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_784
timestamp 1679581782
transform 1 0 75840 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_791
timestamp 1679581782
transform 1 0 76512 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_798
timestamp 1679581782
transform 1 0 77184 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_805
timestamp 1679581782
transform 1 0 77856 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_812
timestamp 1679581782
transform 1 0 78528 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_819
timestamp 1679581782
transform 1 0 79200 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_826
timestamp 1679581782
transform 1 0 79872 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_833
timestamp 1679581782
transform 1 0 80544 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_840
timestamp 1679581782
transform 1 0 81216 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_847
timestamp 1679581782
transform 1 0 81888 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_854
timestamp 1679581782
transform 1 0 82560 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_861
timestamp 1679581782
transform 1 0 83232 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_868
timestamp 1679581782
transform 1 0 83904 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_875
timestamp 1679581782
transform 1 0 84576 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_882
timestamp 1679581782
transform 1 0 85248 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_889
timestamp 1679581782
transform 1 0 85920 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_896
timestamp 1679581782
transform 1 0 86592 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_903
timestamp 1679581782
transform 1 0 87264 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_910
timestamp 1679581782
transform 1 0 87936 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_917
timestamp 1679581782
transform 1 0 88608 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_924
timestamp 1679581782
transform 1 0 89280 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_931
timestamp 1679581782
transform 1 0 89952 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_938
timestamp 1679581782
transform 1 0 90624 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_945
timestamp 1679581782
transform 1 0 91296 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_952
timestamp 1679581782
transform 1 0 91968 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_959
timestamp 1679581782
transform 1 0 92640 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_966
timestamp 1679581782
transform 1 0 93312 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_973
timestamp 1679581782
transform 1 0 93984 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_980
timestamp 1679581782
transform 1 0 94656 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_987
timestamp 1679581782
transform 1 0 95328 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_994
timestamp 1679581782
transform 1 0 96000 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_1001
timestamp 1679581782
transform 1 0 96672 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_1008
timestamp 1679581782
transform 1 0 97344 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_1015
timestamp 1679581782
transform 1 0 98016 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_1022
timestamp 1679581782
transform 1 0 98688 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_4
timestamp 1679581782
transform 1 0 960 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_11
timestamp 1679581782
transform 1 0 1632 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_18
timestamp 1679581782
transform 1 0 2304 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_25
timestamp 1679581782
transform 1 0 2976 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_32
timestamp 1679581782
transform 1 0 3648 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_39
timestamp 1679581782
transform 1 0 4320 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_46
timestamp 1679581782
transform 1 0 4992 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_53
timestamp 1679581782
transform 1 0 5664 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_60
timestamp 1679581782
transform 1 0 6336 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_67
timestamp 1679581782
transform 1 0 7008 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_74
timestamp 1679581782
transform 1 0 7680 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_81
timestamp 1679581782
transform 1 0 8352 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_88
timestamp 1679581782
transform 1 0 9024 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_95
timestamp 1679581782
transform 1 0 9696 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_102
timestamp 1679581782
transform 1 0 10368 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_109
timestamp 1679581782
transform 1 0 11040 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_116
timestamp 1679581782
transform 1 0 11712 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_123
timestamp 1679581782
transform 1 0 12384 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_130
timestamp 1679581782
transform 1 0 13056 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_137
timestamp 1679581782
transform 1 0 13728 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_144
timestamp 1679581782
transform 1 0 14400 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_151
timestamp 1679581782
transform 1 0 15072 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_158
timestamp 1679581782
transform 1 0 15744 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_165
timestamp 1679581782
transform 1 0 16416 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_172
timestamp 1679581782
transform 1 0 17088 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_179
timestamp 1679581782
transform 1 0 17760 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_186
timestamp 1679581782
transform 1 0 18432 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_193
timestamp 1679581782
transform 1 0 19104 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_200
timestamp 1679581782
transform 1 0 19776 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_207
timestamp 1679581782
transform 1 0 20448 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_214
timestamp 1679581782
transform 1 0 21120 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_221
timestamp 1679581782
transform 1 0 21792 0 1 14364
box -48 -56 720 834
use sg13g2_fill_1  FILLER_18_228
timestamp 1677579658
transform 1 0 22464 0 1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_18_256
timestamp 1679581782
transform 1 0 25152 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_263
timestamp 1679581782
transform 1 0 25824 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_270
timestamp 1679581782
transform 1 0 26496 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_277
timestamp 1679581782
transform 1 0 27168 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_284
timestamp 1679581782
transform 1 0 27840 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_291
timestamp 1679581782
transform 1 0 28512 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_298
timestamp 1679581782
transform 1 0 29184 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_305
timestamp 1679581782
transform 1 0 29856 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_312
timestamp 1679581782
transform 1 0 30528 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_319
timestamp 1679581782
transform 1 0 31200 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_326
timestamp 1679581782
transform 1 0 31872 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_333
timestamp 1679581782
transform 1 0 32544 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_340
timestamp 1679581782
transform 1 0 33216 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_347
timestamp 1679581782
transform 1 0 33888 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_354
timestamp 1679581782
transform 1 0 34560 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_361
timestamp 1679581782
transform 1 0 35232 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_368
timestamp 1679581782
transform 1 0 35904 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_375
timestamp 1679581782
transform 1 0 36576 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_382
timestamp 1679581782
transform 1 0 37248 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_389
timestamp 1679581782
transform 1 0 37920 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_396
timestamp 1679581782
transform 1 0 38592 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_403
timestamp 1679581782
transform 1 0 39264 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_410
timestamp 1679581782
transform 1 0 39936 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_417
timestamp 1679581782
transform 1 0 40608 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_424
timestamp 1679581782
transform 1 0 41280 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_431
timestamp 1679581782
transform 1 0 41952 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_438
timestamp 1679581782
transform 1 0 42624 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_445
timestamp 1679581782
transform 1 0 43296 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_452
timestamp 1679581782
transform 1 0 43968 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_459
timestamp 1679581782
transform 1 0 44640 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_466
timestamp 1679581782
transform 1 0 45312 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_473
timestamp 1679581782
transform 1 0 45984 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_480
timestamp 1679581782
transform 1 0 46656 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_487
timestamp 1679581782
transform 1 0 47328 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_494
timestamp 1679581782
transform 1 0 48000 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_501
timestamp 1679581782
transform 1 0 48672 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_508
timestamp 1679581782
transform 1 0 49344 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_515
timestamp 1679581782
transform 1 0 50016 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_522
timestamp 1679581782
transform 1 0 50688 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_529
timestamp 1679581782
transform 1 0 51360 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_536
timestamp 1679581782
transform 1 0 52032 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_543
timestamp 1679581782
transform 1 0 52704 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_550
timestamp 1679581782
transform 1 0 53376 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_557
timestamp 1679581782
transform 1 0 54048 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_564
timestamp 1679581782
transform 1 0 54720 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_571
timestamp 1679581782
transform 1 0 55392 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_578
timestamp 1679581782
transform 1 0 56064 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_585
timestamp 1679581782
transform 1 0 56736 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_592
timestamp 1679581782
transform 1 0 57408 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_599
timestamp 1679581782
transform 1 0 58080 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_606
timestamp 1679581782
transform 1 0 58752 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_613
timestamp 1679581782
transform 1 0 59424 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_620
timestamp 1679581782
transform 1 0 60096 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_627
timestamp 1679581782
transform 1 0 60768 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_634
timestamp 1679581782
transform 1 0 61440 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_641
timestamp 1679581782
transform 1 0 62112 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_648
timestamp 1679581782
transform 1 0 62784 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_655
timestamp 1679581782
transform 1 0 63456 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_662
timestamp 1679581782
transform 1 0 64128 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_669
timestamp 1679581782
transform 1 0 64800 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_676
timestamp 1679581782
transform 1 0 65472 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_683
timestamp 1679581782
transform 1 0 66144 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_690
timestamp 1679581782
transform 1 0 66816 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_697
timestamp 1679581782
transform 1 0 67488 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_704
timestamp 1679581782
transform 1 0 68160 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_711
timestamp 1679581782
transform 1 0 68832 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_718
timestamp 1679581782
transform 1 0 69504 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_725
timestamp 1679581782
transform 1 0 70176 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_732
timestamp 1679581782
transform 1 0 70848 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_739
timestamp 1679581782
transform 1 0 71520 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_746
timestamp 1679581782
transform 1 0 72192 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_753
timestamp 1679581782
transform 1 0 72864 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_760
timestamp 1679581782
transform 1 0 73536 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_767
timestamp 1679581782
transform 1 0 74208 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_774
timestamp 1679581782
transform 1 0 74880 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_781
timestamp 1679581782
transform 1 0 75552 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_788
timestamp 1679581782
transform 1 0 76224 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_795
timestamp 1679581782
transform 1 0 76896 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_802
timestamp 1679581782
transform 1 0 77568 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_809
timestamp 1679581782
transform 1 0 78240 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_816
timestamp 1679581782
transform 1 0 78912 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_823
timestamp 1679581782
transform 1 0 79584 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_830
timestamp 1679581782
transform 1 0 80256 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_837
timestamp 1679581782
transform 1 0 80928 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_844
timestamp 1679581782
transform 1 0 81600 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_851
timestamp 1679581782
transform 1 0 82272 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_858
timestamp 1679581782
transform 1 0 82944 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_865
timestamp 1679581782
transform 1 0 83616 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_872
timestamp 1679581782
transform 1 0 84288 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_879
timestamp 1679581782
transform 1 0 84960 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_886
timestamp 1679581782
transform 1 0 85632 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_893
timestamp 1679581782
transform 1 0 86304 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_900
timestamp 1679581782
transform 1 0 86976 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_907
timestamp 1679581782
transform 1 0 87648 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_914
timestamp 1679581782
transform 1 0 88320 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_921
timestamp 1679581782
transform 1 0 88992 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_928
timestamp 1679581782
transform 1 0 89664 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_935
timestamp 1679581782
transform 1 0 90336 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_942
timestamp 1679581782
transform 1 0 91008 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_949
timestamp 1679581782
transform 1 0 91680 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_956
timestamp 1679581782
transform 1 0 92352 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_963
timestamp 1679581782
transform 1 0 93024 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_970
timestamp 1679581782
transform 1 0 93696 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_977
timestamp 1679581782
transform 1 0 94368 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_984
timestamp 1679581782
transform 1 0 95040 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_991
timestamp 1679581782
transform 1 0 95712 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_998
timestamp 1679581782
transform 1 0 96384 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_1005
timestamp 1679581782
transform 1 0 97056 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_1012
timestamp 1679581782
transform 1 0 97728 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_1019
timestamp 1679581782
transform 1 0 98400 0 1 14364
box -48 -56 720 834
use sg13g2_fill_2  FILLER_18_1026
timestamp 1677580104
transform 1 0 99072 0 1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_18_1028
timestamp 1677579658
transform 1 0 99264 0 1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_19_4
timestamp 1679581782
transform 1 0 960 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_11
timestamp 1679581782
transform 1 0 1632 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_18
timestamp 1679581782
transform 1 0 2304 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_25
timestamp 1679581782
transform 1 0 2976 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_32
timestamp 1679581782
transform 1 0 3648 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_39
timestamp 1679581782
transform 1 0 4320 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_46
timestamp 1679581782
transform 1 0 4992 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_53
timestamp 1679581782
transform 1 0 5664 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_60
timestamp 1679581782
transform 1 0 6336 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_67
timestamp 1679581782
transform 1 0 7008 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_74
timestamp 1679581782
transform 1 0 7680 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_81
timestamp 1679581782
transform 1 0 8352 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_88
timestamp 1679581782
transform 1 0 9024 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_95
timestamp 1679581782
transform 1 0 9696 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_102
timestamp 1679581782
transform 1 0 10368 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_109
timestamp 1679581782
transform 1 0 11040 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_116
timestamp 1679581782
transform 1 0 11712 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_123
timestamp 1679581782
transform 1 0 12384 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_130
timestamp 1679581782
transform 1 0 13056 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_137
timestamp 1679581782
transform 1 0 13728 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_144
timestamp 1679581782
transform 1 0 14400 0 -1 15876
box -48 -56 720 834
use sg13g2_fill_2  FILLER_19_151
timestamp 1677580104
transform 1 0 15072 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_19_153
timestamp 1677579658
transform 1 0 15264 0 -1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_19_181
timestamp 1677580104
transform 1 0 17952 0 -1 15876
box -48 -56 240 834
use sg13g2_decap_8  FILLER_19_192
timestamp 1679581782
transform 1 0 19008 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_199
timestamp 1679581782
transform 1 0 19680 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_206
timestamp 1679581782
transform 1 0 20352 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_213
timestamp 1679581782
transform 1 0 21024 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_220
timestamp 1679581782
transform 1 0 21696 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_227
timestamp 1679581782
transform 1 0 22368 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_234
timestamp 1679581782
transform 1 0 23040 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_241
timestamp 1679581782
transform 1 0 23712 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_248
timestamp 1679581782
transform 1 0 24384 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_255
timestamp 1679581782
transform 1 0 25056 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_262
timestamp 1679581782
transform 1 0 25728 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_269
timestamp 1679581782
transform 1 0 26400 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_276
timestamp 1679581782
transform 1 0 27072 0 -1 15876
box -48 -56 720 834
use sg13g2_fill_1  FILLER_19_283
timestamp 1677579658
transform 1 0 27744 0 -1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_19_290
timestamp 1679581782
transform 1 0 28416 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_297
timestamp 1679581782
transform 1 0 29088 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_304
timestamp 1679581782
transform 1 0 29760 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_311
timestamp 1679581782
transform 1 0 30432 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_318
timestamp 1679581782
transform 1 0 31104 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_325
timestamp 1679581782
transform 1 0 31776 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_332
timestamp 1679581782
transform 1 0 32448 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_339
timestamp 1679581782
transform 1 0 33120 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_346
timestamp 1679581782
transform 1 0 33792 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_353
timestamp 1679581782
transform 1 0 34464 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_360
timestamp 1679581782
transform 1 0 35136 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_367
timestamp 1679581782
transform 1 0 35808 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_374
timestamp 1679581782
transform 1 0 36480 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_4  FILLER_19_381
timestamp 1679577901
transform 1 0 37152 0 -1 15876
box -48 -56 432 834
use sg13g2_decap_8  FILLER_19_412
timestamp 1679581782
transform 1 0 40128 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_419
timestamp 1679581782
transform 1 0 40800 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_426
timestamp 1679581782
transform 1 0 41472 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_433
timestamp 1679581782
transform 1 0 42144 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_440
timestamp 1679581782
transform 1 0 42816 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_447
timestamp 1679581782
transform 1 0 43488 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_454
timestamp 1679581782
transform 1 0 44160 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_461
timestamp 1679581782
transform 1 0 44832 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_468
timestamp 1679581782
transform 1 0 45504 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_475
timestamp 1679581782
transform 1 0 46176 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_482
timestamp 1679581782
transform 1 0 46848 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_489
timestamp 1679581782
transform 1 0 47520 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_496
timestamp 1679581782
transform 1 0 48192 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_503
timestamp 1679581782
transform 1 0 48864 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_510
timestamp 1679581782
transform 1 0 49536 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_517
timestamp 1679581782
transform 1 0 50208 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_524
timestamp 1679581782
transform 1 0 50880 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_531
timestamp 1679581782
transform 1 0 51552 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_538
timestamp 1679581782
transform 1 0 52224 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_545
timestamp 1679581782
transform 1 0 52896 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_552
timestamp 1679581782
transform 1 0 53568 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_559
timestamp 1679581782
transform 1 0 54240 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_566
timestamp 1679581782
transform 1 0 54912 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_573
timestamp 1679581782
transform 1 0 55584 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_580
timestamp 1679581782
transform 1 0 56256 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_587
timestamp 1679581782
transform 1 0 56928 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_594
timestamp 1679581782
transform 1 0 57600 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_601
timestamp 1679581782
transform 1 0 58272 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_608
timestamp 1679581782
transform 1 0 58944 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_615
timestamp 1679581782
transform 1 0 59616 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_622
timestamp 1679581782
transform 1 0 60288 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_629
timestamp 1679581782
transform 1 0 60960 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_636
timestamp 1679581782
transform 1 0 61632 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_643
timestamp 1679581782
transform 1 0 62304 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_650
timestamp 1679581782
transform 1 0 62976 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_657
timestamp 1679581782
transform 1 0 63648 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_664
timestamp 1679581782
transform 1 0 64320 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_671
timestamp 1679581782
transform 1 0 64992 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_678
timestamp 1679581782
transform 1 0 65664 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_685
timestamp 1679581782
transform 1 0 66336 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_692
timestamp 1679581782
transform 1 0 67008 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_699
timestamp 1679581782
transform 1 0 67680 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_706
timestamp 1679581782
transform 1 0 68352 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_713
timestamp 1679581782
transform 1 0 69024 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_720
timestamp 1679581782
transform 1 0 69696 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_727
timestamp 1679581782
transform 1 0 70368 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_734
timestamp 1679581782
transform 1 0 71040 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_741
timestamp 1679581782
transform 1 0 71712 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_748
timestamp 1679581782
transform 1 0 72384 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_755
timestamp 1679581782
transform 1 0 73056 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_762
timestamp 1679581782
transform 1 0 73728 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_769
timestamp 1679581782
transform 1 0 74400 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_776
timestamp 1679581782
transform 1 0 75072 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_783
timestamp 1679581782
transform 1 0 75744 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_790
timestamp 1679581782
transform 1 0 76416 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_797
timestamp 1679581782
transform 1 0 77088 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_804
timestamp 1679581782
transform 1 0 77760 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_811
timestamp 1679581782
transform 1 0 78432 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_818
timestamp 1679581782
transform 1 0 79104 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_825
timestamp 1679581782
transform 1 0 79776 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_832
timestamp 1679581782
transform 1 0 80448 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_839
timestamp 1679581782
transform 1 0 81120 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_846
timestamp 1679581782
transform 1 0 81792 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_853
timestamp 1679581782
transform 1 0 82464 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_860
timestamp 1679581782
transform 1 0 83136 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_867
timestamp 1679581782
transform 1 0 83808 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_874
timestamp 1679581782
transform 1 0 84480 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_881
timestamp 1679581782
transform 1 0 85152 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_888
timestamp 1679581782
transform 1 0 85824 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_895
timestamp 1679581782
transform 1 0 86496 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_902
timestamp 1679581782
transform 1 0 87168 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_909
timestamp 1679581782
transform 1 0 87840 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_916
timestamp 1679581782
transform 1 0 88512 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_923
timestamp 1679581782
transform 1 0 89184 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_930
timestamp 1679581782
transform 1 0 89856 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_937
timestamp 1679581782
transform 1 0 90528 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_944
timestamp 1679581782
transform 1 0 91200 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_951
timestamp 1679581782
transform 1 0 91872 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_958
timestamp 1679581782
transform 1 0 92544 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_965
timestamp 1679581782
transform 1 0 93216 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_972
timestamp 1679581782
transform 1 0 93888 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_979
timestamp 1679581782
transform 1 0 94560 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_986
timestamp 1679581782
transform 1 0 95232 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_993
timestamp 1679581782
transform 1 0 95904 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_1000
timestamp 1679581782
transform 1 0 96576 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_1007
timestamp 1679581782
transform 1 0 97248 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_1014
timestamp 1679581782
transform 1 0 97920 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_1021
timestamp 1679581782
transform 1 0 98592 0 -1 15876
box -48 -56 720 834
use sg13g2_fill_1  FILLER_19_1028
timestamp 1677579658
transform 1 0 99264 0 -1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_20_4
timestamp 1679581782
transform 1 0 960 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_11
timestamp 1679581782
transform 1 0 1632 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_18
timestamp 1679581782
transform 1 0 2304 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_25
timestamp 1679581782
transform 1 0 2976 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_32
timestamp 1679581782
transform 1 0 3648 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_39
timestamp 1679581782
transform 1 0 4320 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_46
timestamp 1679581782
transform 1 0 4992 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_53
timestamp 1679581782
transform 1 0 5664 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_60
timestamp 1679581782
transform 1 0 6336 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_67
timestamp 1679581782
transform 1 0 7008 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_74
timestamp 1679581782
transform 1 0 7680 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_81
timestamp 1679581782
transform 1 0 8352 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_88
timestamp 1679581782
transform 1 0 9024 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_95
timestamp 1679581782
transform 1 0 9696 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_102
timestamp 1679581782
transform 1 0 10368 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_109
timestamp 1679581782
transform 1 0 11040 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_116
timestamp 1679581782
transform 1 0 11712 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_123
timestamp 1679581782
transform 1 0 12384 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_130
timestamp 1679581782
transform 1 0 13056 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_137
timestamp 1679581782
transform 1 0 13728 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_144
timestamp 1679581782
transform 1 0 14400 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_151
timestamp 1679581782
transform 1 0 15072 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_158
timestamp 1679581782
transform 1 0 15744 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_165
timestamp 1679581782
transform 1 0 16416 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_172
timestamp 1679581782
transform 1 0 17088 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_179
timestamp 1679581782
transform 1 0 17760 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_186
timestamp 1679581782
transform 1 0 18432 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_193
timestamp 1679581782
transform 1 0 19104 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_200
timestamp 1679581782
transform 1 0 19776 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_207
timestamp 1679581782
transform 1 0 20448 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_214
timestamp 1679581782
transform 1 0 21120 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_221
timestamp 1679581782
transform 1 0 21792 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_228
timestamp 1679581782
transform 1 0 22464 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_235
timestamp 1679581782
transform 1 0 23136 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_242
timestamp 1679581782
transform 1 0 23808 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_249
timestamp 1679581782
transform 1 0 24480 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_256
timestamp 1679581782
transform 1 0 25152 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_263
timestamp 1679581782
transform 1 0 25824 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_270
timestamp 1679581782
transform 1 0 26496 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_277
timestamp 1679581782
transform 1 0 27168 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_284
timestamp 1679581782
transform 1 0 27840 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_291
timestamp 1679581782
transform 1 0 28512 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_298
timestamp 1679581782
transform 1 0 29184 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_305
timestamp 1679581782
transform 1 0 29856 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_312
timestamp 1679581782
transform 1 0 30528 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_319
timestamp 1679581782
transform 1 0 31200 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_326
timestamp 1679581782
transform 1 0 31872 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_333
timestamp 1679581782
transform 1 0 32544 0 1 15876
box -48 -56 720 834
use sg13g2_decap_4  FILLER_20_340
timestamp 1679577901
transform 1 0 33216 0 1 15876
box -48 -56 432 834
use sg13g2_fill_1  FILLER_20_344
timestamp 1677579658
transform 1 0 33600 0 1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_20_351
timestamp 1679581782
transform 1 0 34272 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_358
timestamp 1679581782
transform 1 0 34944 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_365
timestamp 1679581782
transform 1 0 35616 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_372
timestamp 1679581782
transform 1 0 36288 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_384
timestamp 1679581782
transform 1 0 37440 0 1 15876
box -48 -56 720 834
use sg13g2_decap_4  FILLER_20_391
timestamp 1679577901
transform 1 0 38112 0 1 15876
box -48 -56 432 834
use sg13g2_decap_8  FILLER_20_404
timestamp 1679581782
transform 1 0 39360 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_411
timestamp 1679581782
transform 1 0 40032 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_418
timestamp 1679581782
transform 1 0 40704 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_425
timestamp 1679581782
transform 1 0 41376 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_432
timestamp 1679581782
transform 1 0 42048 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_439
timestamp 1679581782
transform 1 0 42720 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_446
timestamp 1679581782
transform 1 0 43392 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_453
timestamp 1679581782
transform 1 0 44064 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_460
timestamp 1679581782
transform 1 0 44736 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_467
timestamp 1679581782
transform 1 0 45408 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_474
timestamp 1679581782
transform 1 0 46080 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_481
timestamp 1679581782
transform 1 0 46752 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_488
timestamp 1679581782
transform 1 0 47424 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_495
timestamp 1679581782
transform 1 0 48096 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_502
timestamp 1679581782
transform 1 0 48768 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_509
timestamp 1679581782
transform 1 0 49440 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_516
timestamp 1679581782
transform 1 0 50112 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_523
timestamp 1679581782
transform 1 0 50784 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_530
timestamp 1679581782
transform 1 0 51456 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_537
timestamp 1679581782
transform 1 0 52128 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_544
timestamp 1679581782
transform 1 0 52800 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_551
timestamp 1679581782
transform 1 0 53472 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_558
timestamp 1679581782
transform 1 0 54144 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_565
timestamp 1679581782
transform 1 0 54816 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_572
timestamp 1679581782
transform 1 0 55488 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_579
timestamp 1679581782
transform 1 0 56160 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_586
timestamp 1679581782
transform 1 0 56832 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_593
timestamp 1679581782
transform 1 0 57504 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_600
timestamp 1679581782
transform 1 0 58176 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_607
timestamp 1679581782
transform 1 0 58848 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_614
timestamp 1679581782
transform 1 0 59520 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_621
timestamp 1679581782
transform 1 0 60192 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_628
timestamp 1679581782
transform 1 0 60864 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_635
timestamp 1679581782
transform 1 0 61536 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_642
timestamp 1679581782
transform 1 0 62208 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_649
timestamp 1679581782
transform 1 0 62880 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_656
timestamp 1679581782
transform 1 0 63552 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_663
timestamp 1679581782
transform 1 0 64224 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_670
timestamp 1679581782
transform 1 0 64896 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_677
timestamp 1679581782
transform 1 0 65568 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_684
timestamp 1679581782
transform 1 0 66240 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_691
timestamp 1679581782
transform 1 0 66912 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_698
timestamp 1679581782
transform 1 0 67584 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_705
timestamp 1679581782
transform 1 0 68256 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_712
timestamp 1679581782
transform 1 0 68928 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_719
timestamp 1679581782
transform 1 0 69600 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_726
timestamp 1679581782
transform 1 0 70272 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_733
timestamp 1679581782
transform 1 0 70944 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_740
timestamp 1679581782
transform 1 0 71616 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_747
timestamp 1679581782
transform 1 0 72288 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_754
timestamp 1679581782
transform 1 0 72960 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_761
timestamp 1679581782
transform 1 0 73632 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_768
timestamp 1679581782
transform 1 0 74304 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_775
timestamp 1679581782
transform 1 0 74976 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_782
timestamp 1679581782
transform 1 0 75648 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_789
timestamp 1679581782
transform 1 0 76320 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_796
timestamp 1679581782
transform 1 0 76992 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_803
timestamp 1679581782
transform 1 0 77664 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_810
timestamp 1679581782
transform 1 0 78336 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_817
timestamp 1679581782
transform 1 0 79008 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_824
timestamp 1679581782
transform 1 0 79680 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_831
timestamp 1679581782
transform 1 0 80352 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_838
timestamp 1679581782
transform 1 0 81024 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_845
timestamp 1679581782
transform 1 0 81696 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_852
timestamp 1679581782
transform 1 0 82368 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_859
timestamp 1679581782
transform 1 0 83040 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_866
timestamp 1679581782
transform 1 0 83712 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_873
timestamp 1679581782
transform 1 0 84384 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_880
timestamp 1679581782
transform 1 0 85056 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_887
timestamp 1679581782
transform 1 0 85728 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_894
timestamp 1679581782
transform 1 0 86400 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_901
timestamp 1679581782
transform 1 0 87072 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_908
timestamp 1679581782
transform 1 0 87744 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_915
timestamp 1679581782
transform 1 0 88416 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_922
timestamp 1679581782
transform 1 0 89088 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_929
timestamp 1679581782
transform 1 0 89760 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_936
timestamp 1679581782
transform 1 0 90432 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_943
timestamp 1679581782
transform 1 0 91104 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_950
timestamp 1679581782
transform 1 0 91776 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_957
timestamp 1679581782
transform 1 0 92448 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_964
timestamp 1679581782
transform 1 0 93120 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_971
timestamp 1679581782
transform 1 0 93792 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_978
timestamp 1679581782
transform 1 0 94464 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_985
timestamp 1679581782
transform 1 0 95136 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_992
timestamp 1679581782
transform 1 0 95808 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_999
timestamp 1679581782
transform 1 0 96480 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_1006
timestamp 1679581782
transform 1 0 97152 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_1013
timestamp 1679581782
transform 1 0 97824 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_1020
timestamp 1679581782
transform 1 0 98496 0 1 15876
box -48 -56 720 834
use sg13g2_fill_2  FILLER_20_1027
timestamp 1677580104
transform 1 0 99168 0 1 15876
box -48 -56 240 834
use sg13g2_decap_8  FILLER_21_4
timestamp 1679581782
transform 1 0 960 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_11
timestamp 1679581782
transform 1 0 1632 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_18
timestamp 1679581782
transform 1 0 2304 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_25
timestamp 1679581782
transform 1 0 2976 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_32
timestamp 1679581782
transform 1 0 3648 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_39
timestamp 1679581782
transform 1 0 4320 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_46
timestamp 1679581782
transform 1 0 4992 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_53
timestamp 1679581782
transform 1 0 5664 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_60
timestamp 1679581782
transform 1 0 6336 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_67
timestamp 1679581782
transform 1 0 7008 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_74
timestamp 1679581782
transform 1 0 7680 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_81
timestamp 1679581782
transform 1 0 8352 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_88
timestamp 1679581782
transform 1 0 9024 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_95
timestamp 1679581782
transform 1 0 9696 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_102
timestamp 1679581782
transform 1 0 10368 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_109
timestamp 1679581782
transform 1 0 11040 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_116
timestamp 1679581782
transform 1 0 11712 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_123
timestamp 1679581782
transform 1 0 12384 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_130
timestamp 1679581782
transform 1 0 13056 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_137
timestamp 1679581782
transform 1 0 13728 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_144
timestamp 1679581782
transform 1 0 14400 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_151
timestamp 1679581782
transform 1 0 15072 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_162
timestamp 1679581782
transform 1 0 16128 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_169
timestamp 1679581782
transform 1 0 16800 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_176
timestamp 1679581782
transform 1 0 17472 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_183
timestamp 1679581782
transform 1 0 18144 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_190
timestamp 1679581782
transform 1 0 18816 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_197
timestamp 1679581782
transform 1 0 19488 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_204
timestamp 1679581782
transform 1 0 20160 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_211
timestamp 1679581782
transform 1 0 20832 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_4  FILLER_21_218
timestamp 1679577901
transform 1 0 21504 0 -1 17388
box -48 -56 432 834
use sg13g2_fill_1  FILLER_21_222
timestamp 1677579658
transform 1 0 21888 0 -1 17388
box -48 -56 144 834
use sg13g2_decap_8  FILLER_21_228
timestamp 1679581782
transform 1 0 22464 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_235
timestamp 1679581782
transform 1 0 23136 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_242
timestamp 1679581782
transform 1 0 23808 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_249
timestamp 1679581782
transform 1 0 24480 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_256
timestamp 1679581782
transform 1 0 25152 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_263
timestamp 1679581782
transform 1 0 25824 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_270
timestamp 1679581782
transform 1 0 26496 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_277
timestamp 1679581782
transform 1 0 27168 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_284
timestamp 1679581782
transform 1 0 27840 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_291
timestamp 1679581782
transform 1 0 28512 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_298
timestamp 1679581782
transform 1 0 29184 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_305
timestamp 1679581782
transform 1 0 29856 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_312
timestamp 1679581782
transform 1 0 30528 0 -1 17388
box -48 -56 720 834
use sg13g2_fill_1  FILLER_21_319
timestamp 1677579658
transform 1 0 31200 0 -1 17388
box -48 -56 144 834
use sg13g2_decap_8  FILLER_21_353
timestamp 1679581782
transform 1 0 34464 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_360
timestamp 1679581782
transform 1 0 35136 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_367
timestamp 1679581782
transform 1 0 35808 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_374
timestamp 1679581782
transform 1 0 36480 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_381
timestamp 1679581782
transform 1 0 37152 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_388
timestamp 1679581782
transform 1 0 37824 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_395
timestamp 1679581782
transform 1 0 38496 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_402
timestamp 1679581782
transform 1 0 39168 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_409
timestamp 1679581782
transform 1 0 39840 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_416
timestamp 1679581782
transform 1 0 40512 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_423
timestamp 1679581782
transform 1 0 41184 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_430
timestamp 1679581782
transform 1 0 41856 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_437
timestamp 1679581782
transform 1 0 42528 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_444
timestamp 1679581782
transform 1 0 43200 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_451
timestamp 1679581782
transform 1 0 43872 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_458
timestamp 1679581782
transform 1 0 44544 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_465
timestamp 1679581782
transform 1 0 45216 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_472
timestamp 1679581782
transform 1 0 45888 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_479
timestamp 1679581782
transform 1 0 46560 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_486
timestamp 1679581782
transform 1 0 47232 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_493
timestamp 1679581782
transform 1 0 47904 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_500
timestamp 1679581782
transform 1 0 48576 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_507
timestamp 1679581782
transform 1 0 49248 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_514
timestamp 1679581782
transform 1 0 49920 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_521
timestamp 1679581782
transform 1 0 50592 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_528
timestamp 1679581782
transform 1 0 51264 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_535
timestamp 1679581782
transform 1 0 51936 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_542
timestamp 1679581782
transform 1 0 52608 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_549
timestamp 1679581782
transform 1 0 53280 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_556
timestamp 1679581782
transform 1 0 53952 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_563
timestamp 1679581782
transform 1 0 54624 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_570
timestamp 1679581782
transform 1 0 55296 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_577
timestamp 1679581782
transform 1 0 55968 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_584
timestamp 1679581782
transform 1 0 56640 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_591
timestamp 1679581782
transform 1 0 57312 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_598
timestamp 1679581782
transform 1 0 57984 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_605
timestamp 1679581782
transform 1 0 58656 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_612
timestamp 1679581782
transform 1 0 59328 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_619
timestamp 1679581782
transform 1 0 60000 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_626
timestamp 1679581782
transform 1 0 60672 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_633
timestamp 1679581782
transform 1 0 61344 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_640
timestamp 1679581782
transform 1 0 62016 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_647
timestamp 1679581782
transform 1 0 62688 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_654
timestamp 1679581782
transform 1 0 63360 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_661
timestamp 1679581782
transform 1 0 64032 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_668
timestamp 1679581782
transform 1 0 64704 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_675
timestamp 1679581782
transform 1 0 65376 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_682
timestamp 1679581782
transform 1 0 66048 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_689
timestamp 1679581782
transform 1 0 66720 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_696
timestamp 1679581782
transform 1 0 67392 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_703
timestamp 1679581782
transform 1 0 68064 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_710
timestamp 1679581782
transform 1 0 68736 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_717
timestamp 1679581782
transform 1 0 69408 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_724
timestamp 1679581782
transform 1 0 70080 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_731
timestamp 1679581782
transform 1 0 70752 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_738
timestamp 1679581782
transform 1 0 71424 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_745
timestamp 1679581782
transform 1 0 72096 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_752
timestamp 1679581782
transform 1 0 72768 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_759
timestamp 1679581782
transform 1 0 73440 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_766
timestamp 1679581782
transform 1 0 74112 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_773
timestamp 1679581782
transform 1 0 74784 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_780
timestamp 1679581782
transform 1 0 75456 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_787
timestamp 1679581782
transform 1 0 76128 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_794
timestamp 1679581782
transform 1 0 76800 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_801
timestamp 1679581782
transform 1 0 77472 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_808
timestamp 1679581782
transform 1 0 78144 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_815
timestamp 1679581782
transform 1 0 78816 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_822
timestamp 1679581782
transform 1 0 79488 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_829
timestamp 1679581782
transform 1 0 80160 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_836
timestamp 1679581782
transform 1 0 80832 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_843
timestamp 1679581782
transform 1 0 81504 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_850
timestamp 1679581782
transform 1 0 82176 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_857
timestamp 1679581782
transform 1 0 82848 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_864
timestamp 1679581782
transform 1 0 83520 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_871
timestamp 1679581782
transform 1 0 84192 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_878
timestamp 1679581782
transform 1 0 84864 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_885
timestamp 1679581782
transform 1 0 85536 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_892
timestamp 1679581782
transform 1 0 86208 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_899
timestamp 1679581782
transform 1 0 86880 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_906
timestamp 1679581782
transform 1 0 87552 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_913
timestamp 1679581782
transform 1 0 88224 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_920
timestamp 1679581782
transform 1 0 88896 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_927
timestamp 1679581782
transform 1 0 89568 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_934
timestamp 1679581782
transform 1 0 90240 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_941
timestamp 1679581782
transform 1 0 90912 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_948
timestamp 1679581782
transform 1 0 91584 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_955
timestamp 1679581782
transform 1 0 92256 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_962
timestamp 1679581782
transform 1 0 92928 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_969
timestamp 1679581782
transform 1 0 93600 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_976
timestamp 1679581782
transform 1 0 94272 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_983
timestamp 1679581782
transform 1 0 94944 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_990
timestamp 1679581782
transform 1 0 95616 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_997
timestamp 1679581782
transform 1 0 96288 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_1004
timestamp 1679581782
transform 1 0 96960 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_1011
timestamp 1679581782
transform 1 0 97632 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_1018
timestamp 1679581782
transform 1 0 98304 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_4  FILLER_21_1025
timestamp 1679577901
transform 1 0 98976 0 -1 17388
box -48 -56 432 834
use sg13g2_decap_8  FILLER_22_4
timestamp 1679581782
transform 1 0 960 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_11
timestamp 1679581782
transform 1 0 1632 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_18
timestamp 1679581782
transform 1 0 2304 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_25
timestamp 1679581782
transform 1 0 2976 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_32
timestamp 1679581782
transform 1 0 3648 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_39
timestamp 1679581782
transform 1 0 4320 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_46
timestamp 1679581782
transform 1 0 4992 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_53
timestamp 1679581782
transform 1 0 5664 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_60
timestamp 1679581782
transform 1 0 6336 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_67
timestamp 1679581782
transform 1 0 7008 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_74
timestamp 1679581782
transform 1 0 7680 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_81
timestamp 1679581782
transform 1 0 8352 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_88
timestamp 1679581782
transform 1 0 9024 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_95
timestamp 1679581782
transform 1 0 9696 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_102
timestamp 1679581782
transform 1 0 10368 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_109
timestamp 1679581782
transform 1 0 11040 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_116
timestamp 1679581782
transform 1 0 11712 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_123
timestamp 1679581782
transform 1 0 12384 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_130
timestamp 1679581782
transform 1 0 13056 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_137
timestamp 1679581782
transform 1 0 13728 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_144
timestamp 1679581782
transform 1 0 14400 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_151
timestamp 1679581782
transform 1 0 15072 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_166
timestamp 1679581782
transform 1 0 16512 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_173
timestamp 1679581782
transform 1 0 17184 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_180
timestamp 1679581782
transform 1 0 17856 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_187
timestamp 1679581782
transform 1 0 18528 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_194
timestamp 1679581782
transform 1 0 19200 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_201
timestamp 1679581782
transform 1 0 19872 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_208
timestamp 1679581782
transform 1 0 20544 0 1 17388
box -48 -56 720 834
use sg13g2_fill_2  FILLER_22_218
timestamp 1677580104
transform 1 0 21504 0 1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_22_223
timestamp 1677579658
transform 1 0 21984 0 1 17388
box -48 -56 144 834
use sg13g2_decap_8  FILLER_22_233
timestamp 1679581782
transform 1 0 22944 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_240
timestamp 1679581782
transform 1 0 23616 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_247
timestamp 1679581782
transform 1 0 24288 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_254
timestamp 1679581782
transform 1 0 24960 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_261
timestamp 1679581782
transform 1 0 25632 0 1 17388
box -48 -56 720 834
use sg13g2_decap_4  FILLER_22_268
timestamp 1679577901
transform 1 0 26304 0 1 17388
box -48 -56 432 834
use sg13g2_decap_8  FILLER_22_299
timestamp 1679581782
transform 1 0 29280 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_306
timestamp 1679581782
transform 1 0 29952 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_313
timestamp 1679581782
transform 1 0 30624 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_320
timestamp 1679581782
transform 1 0 31296 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_327
timestamp 1679581782
transform 1 0 31968 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_334
timestamp 1679581782
transform 1 0 32640 0 1 17388
box -48 -56 720 834
use sg13g2_fill_2  FILLER_22_341
timestamp 1677580104
transform 1 0 33312 0 1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_22_343
timestamp 1677579658
transform 1 0 33504 0 1 17388
box -48 -56 144 834
use sg13g2_decap_8  FILLER_22_348
timestamp 1679581782
transform 1 0 33984 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_355
timestamp 1679581782
transform 1 0 34656 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_362
timestamp 1679581782
transform 1 0 35328 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_369
timestamp 1679581782
transform 1 0 36000 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_376
timestamp 1679581782
transform 1 0 36672 0 1 17388
box -48 -56 720 834
use sg13g2_decap_4  FILLER_22_383
timestamp 1679577901
transform 1 0 37344 0 1 17388
box -48 -56 432 834
use sg13g2_fill_1  FILLER_22_387
timestamp 1677579658
transform 1 0 37728 0 1 17388
box -48 -56 144 834
use sg13g2_decap_8  FILLER_22_401
timestamp 1679581782
transform 1 0 39072 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_408
timestamp 1679581782
transform 1 0 39744 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_415
timestamp 1679581782
transform 1 0 40416 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_422
timestamp 1679581782
transform 1 0 41088 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_429
timestamp 1679581782
transform 1 0 41760 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_436
timestamp 1679581782
transform 1 0 42432 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_443
timestamp 1679581782
transform 1 0 43104 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_450
timestamp 1679581782
transform 1 0 43776 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_457
timestamp 1679581782
transform 1 0 44448 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_464
timestamp 1679581782
transform 1 0 45120 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_471
timestamp 1679581782
transform 1 0 45792 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_478
timestamp 1679581782
transform 1 0 46464 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_485
timestamp 1679581782
transform 1 0 47136 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_492
timestamp 1679581782
transform 1 0 47808 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_499
timestamp 1679581782
transform 1 0 48480 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_506
timestamp 1679581782
transform 1 0 49152 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_513
timestamp 1679581782
transform 1 0 49824 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_520
timestamp 1679581782
transform 1 0 50496 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_527
timestamp 1679581782
transform 1 0 51168 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_534
timestamp 1679581782
transform 1 0 51840 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_541
timestamp 1679581782
transform 1 0 52512 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_548
timestamp 1679581782
transform 1 0 53184 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_555
timestamp 1679581782
transform 1 0 53856 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_562
timestamp 1679581782
transform 1 0 54528 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_569
timestamp 1679581782
transform 1 0 55200 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_576
timestamp 1679581782
transform 1 0 55872 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_583
timestamp 1679581782
transform 1 0 56544 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_590
timestamp 1679581782
transform 1 0 57216 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_597
timestamp 1679581782
transform 1 0 57888 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_604
timestamp 1679581782
transform 1 0 58560 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_611
timestamp 1679581782
transform 1 0 59232 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_618
timestamp 1679581782
transform 1 0 59904 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_625
timestamp 1679581782
transform 1 0 60576 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_632
timestamp 1679581782
transform 1 0 61248 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_639
timestamp 1679581782
transform 1 0 61920 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_646
timestamp 1679581782
transform 1 0 62592 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_653
timestamp 1679581782
transform 1 0 63264 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_660
timestamp 1679581782
transform 1 0 63936 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_667
timestamp 1679581782
transform 1 0 64608 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_674
timestamp 1679581782
transform 1 0 65280 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_681
timestamp 1679581782
transform 1 0 65952 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_688
timestamp 1679581782
transform 1 0 66624 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_695
timestamp 1679581782
transform 1 0 67296 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_702
timestamp 1679581782
transform 1 0 67968 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_709
timestamp 1679581782
transform 1 0 68640 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_716
timestamp 1679581782
transform 1 0 69312 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_723
timestamp 1679581782
transform 1 0 69984 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_730
timestamp 1679581782
transform 1 0 70656 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_737
timestamp 1679581782
transform 1 0 71328 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_744
timestamp 1679581782
transform 1 0 72000 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_751
timestamp 1679581782
transform 1 0 72672 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_758
timestamp 1679581782
transform 1 0 73344 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_765
timestamp 1679581782
transform 1 0 74016 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_772
timestamp 1679581782
transform 1 0 74688 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_779
timestamp 1679581782
transform 1 0 75360 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_786
timestamp 1679581782
transform 1 0 76032 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_793
timestamp 1679581782
transform 1 0 76704 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_800
timestamp 1679581782
transform 1 0 77376 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_807
timestamp 1679581782
transform 1 0 78048 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_814
timestamp 1679581782
transform 1 0 78720 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_821
timestamp 1679581782
transform 1 0 79392 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_828
timestamp 1679581782
transform 1 0 80064 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_835
timestamp 1679581782
transform 1 0 80736 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_842
timestamp 1679581782
transform 1 0 81408 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_849
timestamp 1679581782
transform 1 0 82080 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_856
timestamp 1679581782
transform 1 0 82752 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_863
timestamp 1679581782
transform 1 0 83424 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_870
timestamp 1679581782
transform 1 0 84096 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_877
timestamp 1679581782
transform 1 0 84768 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_884
timestamp 1679581782
transform 1 0 85440 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_891
timestamp 1679581782
transform 1 0 86112 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_898
timestamp 1679581782
transform 1 0 86784 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_905
timestamp 1679581782
transform 1 0 87456 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_912
timestamp 1679581782
transform 1 0 88128 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_919
timestamp 1679581782
transform 1 0 88800 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_926
timestamp 1679581782
transform 1 0 89472 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_933
timestamp 1679581782
transform 1 0 90144 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_940
timestamp 1679581782
transform 1 0 90816 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_947
timestamp 1679581782
transform 1 0 91488 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_954
timestamp 1679581782
transform 1 0 92160 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_961
timestamp 1679581782
transform 1 0 92832 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_968
timestamp 1679581782
transform 1 0 93504 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_975
timestamp 1679581782
transform 1 0 94176 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_982
timestamp 1679581782
transform 1 0 94848 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_989
timestamp 1679581782
transform 1 0 95520 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_996
timestamp 1679581782
transform 1 0 96192 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_1003
timestamp 1679581782
transform 1 0 96864 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_1010
timestamp 1679581782
transform 1 0 97536 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_1017
timestamp 1679581782
transform 1 0 98208 0 1 17388
box -48 -56 720 834
use sg13g2_decap_4  FILLER_22_1024
timestamp 1679577901
transform 1 0 98880 0 1 17388
box -48 -56 432 834
use sg13g2_fill_1  FILLER_22_1028
timestamp 1677579658
transform 1 0 99264 0 1 17388
box -48 -56 144 834
use sg13g2_decap_8  FILLER_23_4
timestamp 1679581782
transform 1 0 960 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_11
timestamp 1679581782
transform 1 0 1632 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_18
timestamp 1679581782
transform 1 0 2304 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_25
timestamp 1679581782
transform 1 0 2976 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_32
timestamp 1679581782
transform 1 0 3648 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_39
timestamp 1679581782
transform 1 0 4320 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_46
timestamp 1679581782
transform 1 0 4992 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_53
timestamp 1679581782
transform 1 0 5664 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_60
timestamp 1679581782
transform 1 0 6336 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_67
timestamp 1679581782
transform 1 0 7008 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_74
timestamp 1679581782
transform 1 0 7680 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_81
timestamp 1679581782
transform 1 0 8352 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_88
timestamp 1679581782
transform 1 0 9024 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_95
timestamp 1679581782
transform 1 0 9696 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_102
timestamp 1679581782
transform 1 0 10368 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_109
timestamp 1679581782
transform 1 0 11040 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_116
timestamp 1679581782
transform 1 0 11712 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_123
timestamp 1679581782
transform 1 0 12384 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_130
timestamp 1679581782
transform 1 0 13056 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_137
timestamp 1679581782
transform 1 0 13728 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_144
timestamp 1679581782
transform 1 0 14400 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_151
timestamp 1679581782
transform 1 0 15072 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_158
timestamp 1679581782
transform 1 0 15744 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_165
timestamp 1679581782
transform 1 0 16416 0 -1 18900
box -48 -56 720 834
use sg13g2_fill_2  FILLER_23_172
timestamp 1677580104
transform 1 0 17088 0 -1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_23_174
timestamp 1677579658
transform 1 0 17280 0 -1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_23_183
timestamp 1679581782
transform 1 0 18144 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_190
timestamp 1679581782
transform 1 0 18816 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_197
timestamp 1679581782
transform 1 0 19488 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_204
timestamp 1679581782
transform 1 0 20160 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_211
timestamp 1679581782
transform 1 0 20832 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_4  FILLER_23_218
timestamp 1679577901
transform 1 0 21504 0 -1 18900
box -48 -56 432 834
use sg13g2_fill_2  FILLER_23_222
timestamp 1677580104
transform 1 0 21888 0 -1 18900
box -48 -56 240 834
use sg13g2_decap_8  FILLER_23_230
timestamp 1679581782
transform 1 0 22656 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_237
timestamp 1679581782
transform 1 0 23328 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_244
timestamp 1679581782
transform 1 0 24000 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_251
timestamp 1679581782
transform 1 0 24672 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_258
timestamp 1679581782
transform 1 0 25344 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_271
timestamp 1679581782
transform 1 0 26592 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_281
timestamp 1679581782
transform 1 0 27552 0 -1 18900
box -48 -56 720 834
use sg13g2_fill_1  FILLER_23_288
timestamp 1677579658
transform 1 0 28224 0 -1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_23_298
timestamp 1679581782
transform 1 0 29184 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_305
timestamp 1679581782
transform 1 0 29856 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_312
timestamp 1679581782
transform 1 0 30528 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_319
timestamp 1679581782
transform 1 0 31200 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_326
timestamp 1679581782
transform 1 0 31872 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_333
timestamp 1679581782
transform 1 0 32544 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_340
timestamp 1679581782
transform 1 0 33216 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_347
timestamp 1679581782
transform 1 0 33888 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_354
timestamp 1679581782
transform 1 0 34560 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_361
timestamp 1679581782
transform 1 0 35232 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_368
timestamp 1679581782
transform 1 0 35904 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_375
timestamp 1679581782
transform 1 0 36576 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_382
timestamp 1679581782
transform 1 0 37248 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_389
timestamp 1679581782
transform 1 0 37920 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_396
timestamp 1679581782
transform 1 0 38592 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_403
timestamp 1679581782
transform 1 0 39264 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_410
timestamp 1679581782
transform 1 0 39936 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_417
timestamp 1679581782
transform 1 0 40608 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_424
timestamp 1679581782
transform 1 0 41280 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_431
timestamp 1679581782
transform 1 0 41952 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_438
timestamp 1679581782
transform 1 0 42624 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_445
timestamp 1679581782
transform 1 0 43296 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_452
timestamp 1679581782
transform 1 0 43968 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_459
timestamp 1679581782
transform 1 0 44640 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_466
timestamp 1679581782
transform 1 0 45312 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_473
timestamp 1679581782
transform 1 0 45984 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_480
timestamp 1679581782
transform 1 0 46656 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_487
timestamp 1679581782
transform 1 0 47328 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_494
timestamp 1679581782
transform 1 0 48000 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_501
timestamp 1679581782
transform 1 0 48672 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_508
timestamp 1679581782
transform 1 0 49344 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_515
timestamp 1679581782
transform 1 0 50016 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_522
timestamp 1679581782
transform 1 0 50688 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_529
timestamp 1679581782
transform 1 0 51360 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_536
timestamp 1679581782
transform 1 0 52032 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_543
timestamp 1679581782
transform 1 0 52704 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_550
timestamp 1679581782
transform 1 0 53376 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_557
timestamp 1679581782
transform 1 0 54048 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_564
timestamp 1679581782
transform 1 0 54720 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_571
timestamp 1679581782
transform 1 0 55392 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_578
timestamp 1679581782
transform 1 0 56064 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_585
timestamp 1679581782
transform 1 0 56736 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_592
timestamp 1679581782
transform 1 0 57408 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_599
timestamp 1679581782
transform 1 0 58080 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_606
timestamp 1679581782
transform 1 0 58752 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_613
timestamp 1679581782
transform 1 0 59424 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_620
timestamp 1679581782
transform 1 0 60096 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_627
timestamp 1679581782
transform 1 0 60768 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_634
timestamp 1679581782
transform 1 0 61440 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_641
timestamp 1679581782
transform 1 0 62112 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_648
timestamp 1679581782
transform 1 0 62784 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_655
timestamp 1679581782
transform 1 0 63456 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_662
timestamp 1679581782
transform 1 0 64128 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_669
timestamp 1679581782
transform 1 0 64800 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_676
timestamp 1679581782
transform 1 0 65472 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_683
timestamp 1679581782
transform 1 0 66144 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_690
timestamp 1679581782
transform 1 0 66816 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_697
timestamp 1679581782
transform 1 0 67488 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_704
timestamp 1679581782
transform 1 0 68160 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_711
timestamp 1679581782
transform 1 0 68832 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_718
timestamp 1679581782
transform 1 0 69504 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_725
timestamp 1679581782
transform 1 0 70176 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_732
timestamp 1679581782
transform 1 0 70848 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_739
timestamp 1679581782
transform 1 0 71520 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_746
timestamp 1679581782
transform 1 0 72192 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_753
timestamp 1679581782
transform 1 0 72864 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_760
timestamp 1679581782
transform 1 0 73536 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_767
timestamp 1679581782
transform 1 0 74208 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_774
timestamp 1679581782
transform 1 0 74880 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_781
timestamp 1679581782
transform 1 0 75552 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_788
timestamp 1679581782
transform 1 0 76224 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_795
timestamp 1679581782
transform 1 0 76896 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_802
timestamp 1679581782
transform 1 0 77568 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_809
timestamp 1679581782
transform 1 0 78240 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_816
timestamp 1679581782
transform 1 0 78912 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_823
timestamp 1679581782
transform 1 0 79584 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_830
timestamp 1679581782
transform 1 0 80256 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_837
timestamp 1679581782
transform 1 0 80928 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_844
timestamp 1679581782
transform 1 0 81600 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_851
timestamp 1679581782
transform 1 0 82272 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_858
timestamp 1679581782
transform 1 0 82944 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_865
timestamp 1679581782
transform 1 0 83616 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_872
timestamp 1679581782
transform 1 0 84288 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_879
timestamp 1679581782
transform 1 0 84960 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_886
timestamp 1679581782
transform 1 0 85632 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_893
timestamp 1679581782
transform 1 0 86304 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_900
timestamp 1679581782
transform 1 0 86976 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_907
timestamp 1679581782
transform 1 0 87648 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_914
timestamp 1679581782
transform 1 0 88320 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_921
timestamp 1679581782
transform 1 0 88992 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_928
timestamp 1679581782
transform 1 0 89664 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_935
timestamp 1679581782
transform 1 0 90336 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_942
timestamp 1679581782
transform 1 0 91008 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_949
timestamp 1679581782
transform 1 0 91680 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_956
timestamp 1679581782
transform 1 0 92352 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_963
timestamp 1679581782
transform 1 0 93024 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_970
timestamp 1679581782
transform 1 0 93696 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_977
timestamp 1679581782
transform 1 0 94368 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_984
timestamp 1679581782
transform 1 0 95040 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_991
timestamp 1679581782
transform 1 0 95712 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_998
timestamp 1679581782
transform 1 0 96384 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_1005
timestamp 1679581782
transform 1 0 97056 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_1012
timestamp 1679581782
transform 1 0 97728 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_1019
timestamp 1679581782
transform 1 0 98400 0 -1 18900
box -48 -56 720 834
use sg13g2_fill_2  FILLER_23_1026
timestamp 1677580104
transform 1 0 99072 0 -1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_23_1028
timestamp 1677579658
transform 1 0 99264 0 -1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_24_4
timestamp 1679581782
transform 1 0 960 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_11
timestamp 1679581782
transform 1 0 1632 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_18
timestamp 1679581782
transform 1 0 2304 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_25
timestamp 1679581782
transform 1 0 2976 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_32
timestamp 1679581782
transform 1 0 3648 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_39
timestamp 1679581782
transform 1 0 4320 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_46
timestamp 1679581782
transform 1 0 4992 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_53
timestamp 1679581782
transform 1 0 5664 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_60
timestamp 1679581782
transform 1 0 6336 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_67
timestamp 1679581782
transform 1 0 7008 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_74
timestamp 1679581782
transform 1 0 7680 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_81
timestamp 1679581782
transform 1 0 8352 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_88
timestamp 1679581782
transform 1 0 9024 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_95
timestamp 1679581782
transform 1 0 9696 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_102
timestamp 1679581782
transform 1 0 10368 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_109
timestamp 1679581782
transform 1 0 11040 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_116
timestamp 1679581782
transform 1 0 11712 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_123
timestamp 1679581782
transform 1 0 12384 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_130
timestamp 1679581782
transform 1 0 13056 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_137
timestamp 1679581782
transform 1 0 13728 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_144
timestamp 1679581782
transform 1 0 14400 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_151
timestamp 1679581782
transform 1 0 15072 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_158
timestamp 1679581782
transform 1 0 15744 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_165
timestamp 1679581782
transform 1 0 16416 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_172
timestamp 1679581782
transform 1 0 17088 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_179
timestamp 1679581782
transform 1 0 17760 0 1 18900
box -48 -56 720 834
use sg13g2_fill_2  FILLER_24_186
timestamp 1677580104
transform 1 0 18432 0 1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_24_188
timestamp 1677579658
transform 1 0 18624 0 1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_24_201
timestamp 1679581782
transform 1 0 19872 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_208
timestamp 1679581782
transform 1 0 20544 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_215
timestamp 1679581782
transform 1 0 21216 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_222
timestamp 1679581782
transform 1 0 21888 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_229
timestamp 1679581782
transform 1 0 22560 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_236
timestamp 1679581782
transform 1 0 23232 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_243
timestamp 1679581782
transform 1 0 23904 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_250
timestamp 1679581782
transform 1 0 24576 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_257
timestamp 1679581782
transform 1 0 25248 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_264
timestamp 1679581782
transform 1 0 25920 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_271
timestamp 1679581782
transform 1 0 26592 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_278
timestamp 1679581782
transform 1 0 27264 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_285
timestamp 1679581782
transform 1 0 27936 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_292
timestamp 1679581782
transform 1 0 28608 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_299
timestamp 1679581782
transform 1 0 29280 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_306
timestamp 1679581782
transform 1 0 29952 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_313
timestamp 1679581782
transform 1 0 30624 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_320
timestamp 1679581782
transform 1 0 31296 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_327
timestamp 1679581782
transform 1 0 31968 0 1 18900
box -48 -56 720 834
use sg13g2_decap_4  FILLER_24_334
timestamp 1679577901
transform 1 0 32640 0 1 18900
box -48 -56 432 834
use sg13g2_decap_8  FILLER_24_351
timestamp 1679581782
transform 1 0 34272 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_358
timestamp 1679581782
transform 1 0 34944 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_365
timestamp 1679581782
transform 1 0 35616 0 1 18900
box -48 -56 720 834
use sg13g2_decap_4  FILLER_24_372
timestamp 1679577901
transform 1 0 36288 0 1 18900
box -48 -56 432 834
use sg13g2_decap_8  FILLER_24_386
timestamp 1679581782
transform 1 0 37632 0 1 18900
box -48 -56 720 834
use sg13g2_decap_4  FILLER_24_393
timestamp 1679577901
transform 1 0 38304 0 1 18900
box -48 -56 432 834
use sg13g2_decap_8  FILLER_24_424
timestamp 1679581782
transform 1 0 41280 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_431
timestamp 1679581782
transform 1 0 41952 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_438
timestamp 1679581782
transform 1 0 42624 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_445
timestamp 1679581782
transform 1 0 43296 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_452
timestamp 1679581782
transform 1 0 43968 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_459
timestamp 1679581782
transform 1 0 44640 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_466
timestamp 1679581782
transform 1 0 45312 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_473
timestamp 1679581782
transform 1 0 45984 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_480
timestamp 1679581782
transform 1 0 46656 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_487
timestamp 1679581782
transform 1 0 47328 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_494
timestamp 1679581782
transform 1 0 48000 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_501
timestamp 1679581782
transform 1 0 48672 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_508
timestamp 1679581782
transform 1 0 49344 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_515
timestamp 1679581782
transform 1 0 50016 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_522
timestamp 1679581782
transform 1 0 50688 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_529
timestamp 1679581782
transform 1 0 51360 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_536
timestamp 1679581782
transform 1 0 52032 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_543
timestamp 1679581782
transform 1 0 52704 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_550
timestamp 1679581782
transform 1 0 53376 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_557
timestamp 1679581782
transform 1 0 54048 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_564
timestamp 1679581782
transform 1 0 54720 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_571
timestamp 1679581782
transform 1 0 55392 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_578
timestamp 1679581782
transform 1 0 56064 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_585
timestamp 1679581782
transform 1 0 56736 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_592
timestamp 1679581782
transform 1 0 57408 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_599
timestamp 1679581782
transform 1 0 58080 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_606
timestamp 1679581782
transform 1 0 58752 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_613
timestamp 1679581782
transform 1 0 59424 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_620
timestamp 1679581782
transform 1 0 60096 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_627
timestamp 1679581782
transform 1 0 60768 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_634
timestamp 1679581782
transform 1 0 61440 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_641
timestamp 1679581782
transform 1 0 62112 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_648
timestamp 1679581782
transform 1 0 62784 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_655
timestamp 1679581782
transform 1 0 63456 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_662
timestamp 1679581782
transform 1 0 64128 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_669
timestamp 1679581782
transform 1 0 64800 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_676
timestamp 1679581782
transform 1 0 65472 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_683
timestamp 1679581782
transform 1 0 66144 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_690
timestamp 1679581782
transform 1 0 66816 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_697
timestamp 1679581782
transform 1 0 67488 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_704
timestamp 1679581782
transform 1 0 68160 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_711
timestamp 1679581782
transform 1 0 68832 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_718
timestamp 1679581782
transform 1 0 69504 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_725
timestamp 1679581782
transform 1 0 70176 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_732
timestamp 1679581782
transform 1 0 70848 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_739
timestamp 1679581782
transform 1 0 71520 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_746
timestamp 1679581782
transform 1 0 72192 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_753
timestamp 1679581782
transform 1 0 72864 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_760
timestamp 1679581782
transform 1 0 73536 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_767
timestamp 1679581782
transform 1 0 74208 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_774
timestamp 1679581782
transform 1 0 74880 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_781
timestamp 1679581782
transform 1 0 75552 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_788
timestamp 1679581782
transform 1 0 76224 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_795
timestamp 1679581782
transform 1 0 76896 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_802
timestamp 1679581782
transform 1 0 77568 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_809
timestamp 1679581782
transform 1 0 78240 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_816
timestamp 1679581782
transform 1 0 78912 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_823
timestamp 1679581782
transform 1 0 79584 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_830
timestamp 1679581782
transform 1 0 80256 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_837
timestamp 1679581782
transform 1 0 80928 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_844
timestamp 1679581782
transform 1 0 81600 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_851
timestamp 1679581782
transform 1 0 82272 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_858
timestamp 1679581782
transform 1 0 82944 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_865
timestamp 1679581782
transform 1 0 83616 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_872
timestamp 1679581782
transform 1 0 84288 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_879
timestamp 1679581782
transform 1 0 84960 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_886
timestamp 1679581782
transform 1 0 85632 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_893
timestamp 1679581782
transform 1 0 86304 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_900
timestamp 1679581782
transform 1 0 86976 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_907
timestamp 1679581782
transform 1 0 87648 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_914
timestamp 1679581782
transform 1 0 88320 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_921
timestamp 1679581782
transform 1 0 88992 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_928
timestamp 1679581782
transform 1 0 89664 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_935
timestamp 1679581782
transform 1 0 90336 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_942
timestamp 1679581782
transform 1 0 91008 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_949
timestamp 1679581782
transform 1 0 91680 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_956
timestamp 1679581782
transform 1 0 92352 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_963
timestamp 1679581782
transform 1 0 93024 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_970
timestamp 1679581782
transform 1 0 93696 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_977
timestamp 1679581782
transform 1 0 94368 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_984
timestamp 1679581782
transform 1 0 95040 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_991
timestamp 1679581782
transform 1 0 95712 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_998
timestamp 1679581782
transform 1 0 96384 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_1005
timestamp 1679581782
transform 1 0 97056 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_1012
timestamp 1679581782
transform 1 0 97728 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_1019
timestamp 1679581782
transform 1 0 98400 0 1 18900
box -48 -56 720 834
use sg13g2_fill_2  FILLER_24_1026
timestamp 1677580104
transform 1 0 99072 0 1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_24_1028
timestamp 1677579658
transform 1 0 99264 0 1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_25_4
timestamp 1679581782
transform 1 0 960 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_11
timestamp 1679581782
transform 1 0 1632 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_18
timestamp 1679581782
transform 1 0 2304 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_25
timestamp 1679581782
transform 1 0 2976 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_32
timestamp 1679581782
transform 1 0 3648 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_39
timestamp 1679581782
transform 1 0 4320 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_46
timestamp 1679581782
transform 1 0 4992 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_53
timestamp 1679581782
transform 1 0 5664 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_60
timestamp 1679581782
transform 1 0 6336 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_67
timestamp 1679581782
transform 1 0 7008 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_74
timestamp 1679581782
transform 1 0 7680 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_81
timestamp 1679581782
transform 1 0 8352 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_88
timestamp 1679581782
transform 1 0 9024 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_95
timestamp 1679581782
transform 1 0 9696 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_102
timestamp 1679581782
transform 1 0 10368 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_109
timestamp 1679581782
transform 1 0 11040 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_116
timestamp 1679581782
transform 1 0 11712 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_123
timestamp 1679581782
transform 1 0 12384 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_130
timestamp 1679581782
transform 1 0 13056 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_137
timestamp 1679581782
transform 1 0 13728 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_144
timestamp 1679581782
transform 1 0 14400 0 -1 20412
box -48 -56 720 834
use sg13g2_fill_2  FILLER_25_151
timestamp 1677580104
transform 1 0 15072 0 -1 20412
box -48 -56 240 834
use sg13g2_decap_8  FILLER_25_161
timestamp 1679581782
transform 1 0 16032 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_168
timestamp 1679581782
transform 1 0 16704 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_175
timestamp 1679581782
transform 1 0 17376 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_182
timestamp 1679581782
transform 1 0 18048 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_189
timestamp 1679581782
transform 1 0 18720 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_196
timestamp 1679581782
transform 1 0 19392 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_203
timestamp 1679581782
transform 1 0 20064 0 -1 20412
box -48 -56 720 834
use sg13g2_fill_2  FILLER_25_210
timestamp 1677580104
transform 1 0 20736 0 -1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_25_212
timestamp 1677579658
transform 1 0 20928 0 -1 20412
box -48 -56 144 834
use sg13g2_fill_2  FILLER_25_218
timestamp 1677580104
transform 1 0 21504 0 -1 20412
box -48 -56 240 834
use sg13g2_decap_4  FILLER_25_225
timestamp 1679577901
transform 1 0 22176 0 -1 20412
box -48 -56 432 834
use sg13g2_fill_2  FILLER_25_229
timestamp 1677580104
transform 1 0 22560 0 -1 20412
box -48 -56 240 834
use sg13g2_decap_8  FILLER_25_248
timestamp 1679581782
transform 1 0 24384 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_255
timestamp 1679581782
transform 1 0 25056 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_262
timestamp 1679581782
transform 1 0 25728 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_269
timestamp 1679581782
transform 1 0 26400 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_276
timestamp 1679581782
transform 1 0 27072 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_283
timestamp 1679581782
transform 1 0 27744 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_290
timestamp 1679581782
transform 1 0 28416 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_297
timestamp 1679581782
transform 1 0 29088 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_304
timestamp 1679581782
transform 1 0 29760 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_311
timestamp 1679581782
transform 1 0 30432 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_318
timestamp 1679581782
transform 1 0 31104 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_325
timestamp 1679581782
transform 1 0 31776 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_332
timestamp 1679581782
transform 1 0 32448 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_339
timestamp 1679581782
transform 1 0 33120 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_346
timestamp 1679581782
transform 1 0 33792 0 -1 20412
box -48 -56 720 834
use sg13g2_fill_2  FILLER_25_353
timestamp 1677580104
transform 1 0 34464 0 -1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_25_355
timestamp 1677579658
transform 1 0 34656 0 -1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_25_360
timestamp 1679581782
transform 1 0 35136 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_367
timestamp 1679581782
transform 1 0 35808 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_374
timestamp 1679581782
transform 1 0 36480 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_381
timestamp 1679581782
transform 1 0 37152 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_388
timestamp 1679581782
transform 1 0 37824 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_395
timestamp 1679581782
transform 1 0 38496 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_411
timestamp 1679581782
transform 1 0 40032 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_418
timestamp 1679581782
transform 1 0 40704 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_425
timestamp 1679581782
transform 1 0 41376 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_432
timestamp 1679581782
transform 1 0 42048 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_439
timestamp 1679581782
transform 1 0 42720 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_446
timestamp 1679581782
transform 1 0 43392 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_453
timestamp 1679581782
transform 1 0 44064 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_460
timestamp 1679581782
transform 1 0 44736 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_467
timestamp 1679581782
transform 1 0 45408 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_474
timestamp 1679581782
transform 1 0 46080 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_481
timestamp 1679581782
transform 1 0 46752 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_488
timestamp 1679581782
transform 1 0 47424 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_495
timestamp 1679581782
transform 1 0 48096 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_502
timestamp 1679581782
transform 1 0 48768 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_509
timestamp 1679581782
transform 1 0 49440 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_516
timestamp 1679581782
transform 1 0 50112 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_523
timestamp 1679581782
transform 1 0 50784 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_530
timestamp 1679581782
transform 1 0 51456 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_537
timestamp 1679581782
transform 1 0 52128 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_544
timestamp 1679581782
transform 1 0 52800 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_551
timestamp 1679581782
transform 1 0 53472 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_558
timestamp 1679581782
transform 1 0 54144 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_565
timestamp 1679581782
transform 1 0 54816 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_572
timestamp 1679581782
transform 1 0 55488 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_579
timestamp 1679581782
transform 1 0 56160 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_586
timestamp 1679581782
transform 1 0 56832 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_593
timestamp 1679581782
transform 1 0 57504 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_600
timestamp 1679581782
transform 1 0 58176 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_607
timestamp 1679581782
transform 1 0 58848 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_614
timestamp 1679581782
transform 1 0 59520 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_621
timestamp 1679581782
transform 1 0 60192 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_628
timestamp 1679581782
transform 1 0 60864 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_635
timestamp 1679581782
transform 1 0 61536 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_642
timestamp 1679581782
transform 1 0 62208 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_649
timestamp 1679581782
transform 1 0 62880 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_656
timestamp 1679581782
transform 1 0 63552 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_663
timestamp 1679581782
transform 1 0 64224 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_670
timestamp 1679581782
transform 1 0 64896 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_677
timestamp 1679581782
transform 1 0 65568 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_684
timestamp 1679581782
transform 1 0 66240 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_691
timestamp 1679581782
transform 1 0 66912 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_698
timestamp 1679581782
transform 1 0 67584 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_705
timestamp 1679581782
transform 1 0 68256 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_712
timestamp 1679581782
transform 1 0 68928 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_719
timestamp 1679581782
transform 1 0 69600 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_726
timestamp 1679581782
transform 1 0 70272 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_733
timestamp 1679581782
transform 1 0 70944 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_740
timestamp 1679581782
transform 1 0 71616 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_747
timestamp 1679581782
transform 1 0 72288 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_754
timestamp 1679581782
transform 1 0 72960 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_761
timestamp 1679581782
transform 1 0 73632 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_768
timestamp 1679581782
transform 1 0 74304 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_775
timestamp 1679581782
transform 1 0 74976 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_782
timestamp 1679581782
transform 1 0 75648 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_789
timestamp 1679581782
transform 1 0 76320 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_796
timestamp 1679581782
transform 1 0 76992 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_803
timestamp 1679581782
transform 1 0 77664 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_810
timestamp 1679581782
transform 1 0 78336 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_817
timestamp 1679581782
transform 1 0 79008 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_824
timestamp 1679581782
transform 1 0 79680 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_831
timestamp 1679581782
transform 1 0 80352 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_838
timestamp 1679581782
transform 1 0 81024 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_845
timestamp 1679581782
transform 1 0 81696 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_852
timestamp 1679581782
transform 1 0 82368 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_859
timestamp 1679581782
transform 1 0 83040 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_866
timestamp 1679581782
transform 1 0 83712 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_873
timestamp 1679581782
transform 1 0 84384 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_880
timestamp 1679581782
transform 1 0 85056 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_887
timestamp 1679581782
transform 1 0 85728 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_894
timestamp 1679581782
transform 1 0 86400 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_901
timestamp 1679581782
transform 1 0 87072 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_908
timestamp 1679581782
transform 1 0 87744 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_915
timestamp 1679581782
transform 1 0 88416 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_922
timestamp 1679581782
transform 1 0 89088 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_929
timestamp 1679581782
transform 1 0 89760 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_936
timestamp 1679581782
transform 1 0 90432 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_943
timestamp 1679581782
transform 1 0 91104 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_950
timestamp 1679581782
transform 1 0 91776 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_957
timestamp 1679581782
transform 1 0 92448 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_964
timestamp 1679581782
transform 1 0 93120 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_971
timestamp 1679581782
transform 1 0 93792 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_978
timestamp 1679581782
transform 1 0 94464 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_985
timestamp 1679581782
transform 1 0 95136 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_992
timestamp 1679581782
transform 1 0 95808 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_999
timestamp 1679581782
transform 1 0 96480 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_1006
timestamp 1679581782
transform 1 0 97152 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_1013
timestamp 1679581782
transform 1 0 97824 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_1020
timestamp 1679581782
transform 1 0 98496 0 -1 20412
box -48 -56 720 834
use sg13g2_fill_2  FILLER_25_1027
timestamp 1677580104
transform 1 0 99168 0 -1 20412
box -48 -56 240 834
use sg13g2_decap_8  FILLER_26_4
timestamp 1679581782
transform 1 0 960 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_11
timestamp 1679581782
transform 1 0 1632 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_18
timestamp 1679581782
transform 1 0 2304 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_25
timestamp 1679581782
transform 1 0 2976 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_32
timestamp 1679581782
transform 1 0 3648 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_39
timestamp 1679581782
transform 1 0 4320 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_46
timestamp 1679581782
transform 1 0 4992 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_53
timestamp 1679581782
transform 1 0 5664 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_60
timestamp 1679581782
transform 1 0 6336 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_67
timestamp 1679581782
transform 1 0 7008 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_74
timestamp 1679581782
transform 1 0 7680 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_81
timestamp 1679581782
transform 1 0 8352 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_88
timestamp 1679581782
transform 1 0 9024 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_95
timestamp 1679581782
transform 1 0 9696 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_102
timestamp 1679581782
transform 1 0 10368 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_109
timestamp 1679581782
transform 1 0 11040 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_116
timestamp 1679581782
transform 1 0 11712 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_123
timestamp 1679581782
transform 1 0 12384 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_130
timestamp 1679581782
transform 1 0 13056 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_137
timestamp 1679581782
transform 1 0 13728 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_144
timestamp 1679581782
transform 1 0 14400 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_151
timestamp 1679581782
transform 1 0 15072 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_158
timestamp 1679581782
transform 1 0 15744 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_165
timestamp 1679581782
transform 1 0 16416 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_172
timestamp 1679581782
transform 1 0 17088 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_179
timestamp 1679581782
transform 1 0 17760 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_186
timestamp 1679581782
transform 1 0 18432 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_200
timestamp 1679581782
transform 1 0 19776 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_207
timestamp 1679581782
transform 1 0 20448 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_214
timestamp 1679581782
transform 1 0 21120 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_221
timestamp 1679581782
transform 1 0 21792 0 1 20412
box -48 -56 720 834
use sg13g2_fill_1  FILLER_26_228
timestamp 1677579658
transform 1 0 22464 0 1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_26_239
timestamp 1679581782
transform 1 0 23520 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_246
timestamp 1679581782
transform 1 0 24192 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_253
timestamp 1679581782
transform 1 0 24864 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_260
timestamp 1679581782
transform 1 0 25536 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_267
timestamp 1679581782
transform 1 0 26208 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_274
timestamp 1679581782
transform 1 0 26880 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_281
timestamp 1679581782
transform 1 0 27552 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_288
timestamp 1679581782
transform 1 0 28224 0 1 20412
box -48 -56 720 834
use sg13g2_fill_2  FILLER_26_295
timestamp 1677580104
transform 1 0 28896 0 1 20412
box -48 -56 240 834
use sg13g2_decap_4  FILLER_26_304
timestamp 1679577901
transform 1 0 29760 0 1 20412
box -48 -56 432 834
use sg13g2_fill_1  FILLER_26_308
timestamp 1677579658
transform 1 0 30144 0 1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_26_322
timestamp 1679581782
transform 1 0 31488 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_329
timestamp 1679581782
transform 1 0 32160 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_336
timestamp 1679581782
transform 1 0 32832 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_343
timestamp 1679581782
transform 1 0 33504 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_350
timestamp 1679581782
transform 1 0 34176 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_357
timestamp 1679581782
transform 1 0 34848 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_364
timestamp 1679581782
transform 1 0 35520 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_371
timestamp 1679581782
transform 1 0 36192 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_378
timestamp 1679581782
transform 1 0 36864 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_385
timestamp 1679581782
transform 1 0 37536 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_392
timestamp 1679581782
transform 1 0 38208 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_399
timestamp 1679581782
transform 1 0 38880 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_406
timestamp 1679581782
transform 1 0 39552 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_413
timestamp 1679581782
transform 1 0 40224 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_420
timestamp 1679581782
transform 1 0 40896 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_427
timestamp 1679581782
transform 1 0 41568 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_434
timestamp 1679581782
transform 1 0 42240 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_441
timestamp 1679581782
transform 1 0 42912 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_448
timestamp 1679581782
transform 1 0 43584 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_455
timestamp 1679581782
transform 1 0 44256 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_462
timestamp 1679581782
transform 1 0 44928 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_469
timestamp 1679581782
transform 1 0 45600 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_476
timestamp 1679581782
transform 1 0 46272 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_483
timestamp 1679581782
transform 1 0 46944 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_490
timestamp 1679581782
transform 1 0 47616 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_497
timestamp 1679581782
transform 1 0 48288 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_504
timestamp 1679581782
transform 1 0 48960 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_511
timestamp 1679581782
transform 1 0 49632 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_518
timestamp 1679581782
transform 1 0 50304 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_525
timestamp 1679581782
transform 1 0 50976 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_532
timestamp 1679581782
transform 1 0 51648 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_539
timestamp 1679581782
transform 1 0 52320 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_546
timestamp 1679581782
transform 1 0 52992 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_553
timestamp 1679581782
transform 1 0 53664 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_560
timestamp 1679581782
transform 1 0 54336 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_567
timestamp 1679581782
transform 1 0 55008 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_574
timestamp 1679581782
transform 1 0 55680 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_581
timestamp 1679581782
transform 1 0 56352 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_588
timestamp 1679581782
transform 1 0 57024 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_595
timestamp 1679581782
transform 1 0 57696 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_602
timestamp 1679581782
transform 1 0 58368 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_609
timestamp 1679581782
transform 1 0 59040 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_616
timestamp 1679581782
transform 1 0 59712 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_623
timestamp 1679581782
transform 1 0 60384 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_630
timestamp 1679581782
transform 1 0 61056 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_637
timestamp 1679581782
transform 1 0 61728 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_644
timestamp 1679581782
transform 1 0 62400 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_651
timestamp 1679581782
transform 1 0 63072 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_658
timestamp 1679581782
transform 1 0 63744 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_665
timestamp 1679581782
transform 1 0 64416 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_672
timestamp 1679581782
transform 1 0 65088 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_679
timestamp 1679581782
transform 1 0 65760 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_686
timestamp 1679581782
transform 1 0 66432 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_693
timestamp 1679581782
transform 1 0 67104 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_700
timestamp 1679581782
transform 1 0 67776 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_707
timestamp 1679581782
transform 1 0 68448 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_714
timestamp 1679581782
transform 1 0 69120 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_721
timestamp 1679581782
transform 1 0 69792 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_728
timestamp 1679581782
transform 1 0 70464 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_735
timestamp 1679581782
transform 1 0 71136 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_742
timestamp 1679581782
transform 1 0 71808 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_749
timestamp 1679581782
transform 1 0 72480 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_756
timestamp 1679581782
transform 1 0 73152 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_763
timestamp 1679581782
transform 1 0 73824 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_770
timestamp 1679581782
transform 1 0 74496 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_777
timestamp 1679581782
transform 1 0 75168 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_784
timestamp 1679581782
transform 1 0 75840 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_791
timestamp 1679581782
transform 1 0 76512 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_798
timestamp 1679581782
transform 1 0 77184 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_805
timestamp 1679581782
transform 1 0 77856 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_812
timestamp 1679581782
transform 1 0 78528 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_819
timestamp 1679581782
transform 1 0 79200 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_826
timestamp 1679581782
transform 1 0 79872 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_833
timestamp 1679581782
transform 1 0 80544 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_840
timestamp 1679581782
transform 1 0 81216 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_847
timestamp 1679581782
transform 1 0 81888 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_854
timestamp 1679581782
transform 1 0 82560 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_861
timestamp 1679581782
transform 1 0 83232 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_868
timestamp 1679581782
transform 1 0 83904 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_875
timestamp 1679581782
transform 1 0 84576 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_882
timestamp 1679581782
transform 1 0 85248 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_889
timestamp 1679581782
transform 1 0 85920 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_896
timestamp 1679581782
transform 1 0 86592 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_903
timestamp 1679581782
transform 1 0 87264 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_910
timestamp 1679581782
transform 1 0 87936 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_917
timestamp 1679581782
transform 1 0 88608 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_924
timestamp 1679581782
transform 1 0 89280 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_931
timestamp 1679581782
transform 1 0 89952 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_938
timestamp 1679581782
transform 1 0 90624 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_945
timestamp 1679581782
transform 1 0 91296 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_952
timestamp 1679581782
transform 1 0 91968 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_959
timestamp 1679581782
transform 1 0 92640 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_966
timestamp 1679581782
transform 1 0 93312 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_973
timestamp 1679581782
transform 1 0 93984 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_980
timestamp 1679581782
transform 1 0 94656 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_987
timestamp 1679581782
transform 1 0 95328 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_994
timestamp 1679581782
transform 1 0 96000 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_1001
timestamp 1679581782
transform 1 0 96672 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_1008
timestamp 1679581782
transform 1 0 97344 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_1015
timestamp 1679581782
transform 1 0 98016 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_1022
timestamp 1679581782
transform 1 0 98688 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_0
timestamp 1679581782
transform 1 0 576 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_7
timestamp 1679581782
transform 1 0 1248 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_14
timestamp 1679581782
transform 1 0 1920 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_21
timestamp 1679581782
transform 1 0 2592 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_28
timestamp 1679581782
transform 1 0 3264 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_35
timestamp 1679581782
transform 1 0 3936 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_42
timestamp 1679581782
transform 1 0 4608 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_49
timestamp 1679581782
transform 1 0 5280 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_56
timestamp 1679581782
transform 1 0 5952 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_63
timestamp 1679581782
transform 1 0 6624 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_70
timestamp 1679581782
transform 1 0 7296 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_77
timestamp 1679581782
transform 1 0 7968 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_84
timestamp 1679581782
transform 1 0 8640 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_91
timestamp 1679581782
transform 1 0 9312 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_98
timestamp 1679581782
transform 1 0 9984 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_105
timestamp 1679581782
transform 1 0 10656 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_112
timestamp 1679581782
transform 1 0 11328 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_119
timestamp 1679581782
transform 1 0 12000 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_126
timestamp 1679581782
transform 1 0 12672 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_133
timestamp 1679581782
transform 1 0 13344 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_140
timestamp 1679581782
transform 1 0 14016 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_147
timestamp 1679581782
transform 1 0 14688 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_154
timestamp 1679581782
transform 1 0 15360 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_161
timestamp 1679581782
transform 1 0 16032 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_168
timestamp 1679581782
transform 1 0 16704 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_175
timestamp 1679581782
transform 1 0 17376 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_182
timestamp 1679581782
transform 1 0 18048 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_189
timestamp 1679581782
transform 1 0 18720 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_196
timestamp 1679581782
transform 1 0 19392 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_203
timestamp 1679581782
transform 1 0 20064 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_210
timestamp 1679581782
transform 1 0 20736 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_217
timestamp 1679581782
transform 1 0 21408 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_224
timestamp 1679581782
transform 1 0 22080 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_231
timestamp 1679581782
transform 1 0 22752 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_238
timestamp 1679581782
transform 1 0 23424 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_245
timestamp 1679581782
transform 1 0 24096 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_252
timestamp 1679581782
transform 1 0 24768 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_259
timestamp 1679581782
transform 1 0 25440 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_266
timestamp 1679581782
transform 1 0 26112 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_273
timestamp 1679581782
transform 1 0 26784 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_280
timestamp 1679581782
transform 1 0 27456 0 -1 21924
box -48 -56 720 834
use sg13g2_fill_1  FILLER_27_287
timestamp 1677579658
transform 1 0 28128 0 -1 21924
box -48 -56 144 834
use sg13g2_decap_8  FILLER_27_301
timestamp 1679581782
transform 1 0 29472 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_308
timestamp 1679581782
transform 1 0 30144 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_315
timestamp 1679581782
transform 1 0 30816 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_322
timestamp 1679581782
transform 1 0 31488 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_329
timestamp 1679581782
transform 1 0 32160 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_336
timestamp 1679581782
transform 1 0 32832 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_343
timestamp 1679581782
transform 1 0 33504 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_350
timestamp 1679581782
transform 1 0 34176 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_357
timestamp 1679581782
transform 1 0 34848 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_364
timestamp 1679581782
transform 1 0 35520 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_371
timestamp 1679581782
transform 1 0 36192 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_378
timestamp 1679581782
transform 1 0 36864 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_385
timestamp 1679581782
transform 1 0 37536 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_392
timestamp 1679581782
transform 1 0 38208 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_399
timestamp 1679581782
transform 1 0 38880 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_406
timestamp 1679581782
transform 1 0 39552 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_413
timestamp 1679581782
transform 1 0 40224 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_420
timestamp 1679581782
transform 1 0 40896 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_427
timestamp 1679581782
transform 1 0 41568 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_434
timestamp 1679581782
transform 1 0 42240 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_441
timestamp 1679581782
transform 1 0 42912 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_448
timestamp 1679581782
transform 1 0 43584 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_455
timestamp 1679581782
transform 1 0 44256 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_462
timestamp 1679581782
transform 1 0 44928 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_469
timestamp 1679581782
transform 1 0 45600 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_476
timestamp 1679581782
transform 1 0 46272 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_483
timestamp 1679581782
transform 1 0 46944 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_490
timestamp 1679581782
transform 1 0 47616 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_497
timestamp 1679581782
transform 1 0 48288 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_504
timestamp 1679581782
transform 1 0 48960 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_511
timestamp 1679581782
transform 1 0 49632 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_518
timestamp 1679581782
transform 1 0 50304 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_525
timestamp 1679581782
transform 1 0 50976 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_532
timestamp 1679581782
transform 1 0 51648 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_539
timestamp 1679581782
transform 1 0 52320 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_546
timestamp 1679581782
transform 1 0 52992 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_553
timestamp 1679581782
transform 1 0 53664 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_560
timestamp 1679581782
transform 1 0 54336 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_567
timestamp 1679581782
transform 1 0 55008 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_574
timestamp 1679581782
transform 1 0 55680 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_581
timestamp 1679581782
transform 1 0 56352 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_588
timestamp 1679581782
transform 1 0 57024 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_595
timestamp 1679581782
transform 1 0 57696 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_602
timestamp 1679581782
transform 1 0 58368 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_609
timestamp 1679581782
transform 1 0 59040 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_616
timestamp 1679581782
transform 1 0 59712 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_623
timestamp 1679581782
transform 1 0 60384 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_630
timestamp 1679581782
transform 1 0 61056 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_637
timestamp 1679581782
transform 1 0 61728 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_644
timestamp 1679581782
transform 1 0 62400 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_651
timestamp 1679581782
transform 1 0 63072 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_658
timestamp 1679581782
transform 1 0 63744 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_665
timestamp 1679581782
transform 1 0 64416 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_672
timestamp 1679581782
transform 1 0 65088 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_679
timestamp 1679581782
transform 1 0 65760 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_686
timestamp 1679581782
transform 1 0 66432 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_693
timestamp 1679581782
transform 1 0 67104 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_700
timestamp 1679581782
transform 1 0 67776 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_707
timestamp 1679581782
transform 1 0 68448 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_714
timestamp 1679581782
transform 1 0 69120 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_721
timestamp 1679581782
transform 1 0 69792 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_728
timestamp 1679581782
transform 1 0 70464 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_735
timestamp 1679581782
transform 1 0 71136 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_742
timestamp 1679581782
transform 1 0 71808 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_749
timestamp 1679581782
transform 1 0 72480 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_756
timestamp 1679581782
transform 1 0 73152 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_763
timestamp 1679581782
transform 1 0 73824 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_770
timestamp 1679581782
transform 1 0 74496 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_777
timestamp 1679581782
transform 1 0 75168 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_784
timestamp 1679581782
transform 1 0 75840 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_791
timestamp 1679581782
transform 1 0 76512 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_798
timestamp 1679581782
transform 1 0 77184 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_805
timestamp 1679581782
transform 1 0 77856 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_812
timestamp 1679581782
transform 1 0 78528 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_819
timestamp 1679581782
transform 1 0 79200 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_826
timestamp 1679581782
transform 1 0 79872 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_833
timestamp 1679581782
transform 1 0 80544 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_840
timestamp 1679581782
transform 1 0 81216 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_847
timestamp 1679581782
transform 1 0 81888 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_854
timestamp 1679581782
transform 1 0 82560 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_861
timestamp 1679581782
transform 1 0 83232 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_868
timestamp 1679581782
transform 1 0 83904 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_875
timestamp 1679581782
transform 1 0 84576 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_882
timestamp 1679581782
transform 1 0 85248 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_889
timestamp 1679581782
transform 1 0 85920 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_896
timestamp 1679581782
transform 1 0 86592 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_903
timestamp 1679581782
transform 1 0 87264 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_910
timestamp 1679581782
transform 1 0 87936 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_917
timestamp 1679581782
transform 1 0 88608 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_924
timestamp 1679581782
transform 1 0 89280 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_931
timestamp 1679581782
transform 1 0 89952 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_938
timestamp 1679581782
transform 1 0 90624 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_945
timestamp 1679581782
transform 1 0 91296 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_952
timestamp 1679581782
transform 1 0 91968 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_959
timestamp 1679581782
transform 1 0 92640 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_966
timestamp 1679581782
transform 1 0 93312 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_973
timestamp 1679581782
transform 1 0 93984 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_980
timestamp 1679581782
transform 1 0 94656 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_987
timestamp 1679581782
transform 1 0 95328 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_994
timestamp 1679581782
transform 1 0 96000 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_1001
timestamp 1679581782
transform 1 0 96672 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_1008
timestamp 1679581782
transform 1 0 97344 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_1015
timestamp 1679581782
transform 1 0 98016 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_1022
timestamp 1679581782
transform 1 0 98688 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_4
timestamp 1679581782
transform 1 0 960 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_11
timestamp 1679581782
transform 1 0 1632 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_18
timestamp 1679581782
transform 1 0 2304 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_25
timestamp 1679581782
transform 1 0 2976 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_32
timestamp 1679581782
transform 1 0 3648 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_39
timestamp 1679581782
transform 1 0 4320 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_46
timestamp 1679581782
transform 1 0 4992 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_53
timestamp 1679581782
transform 1 0 5664 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_60
timestamp 1679581782
transform 1 0 6336 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_67
timestamp 1679581782
transform 1 0 7008 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_74
timestamp 1679581782
transform 1 0 7680 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_81
timestamp 1679581782
transform 1 0 8352 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_88
timestamp 1679581782
transform 1 0 9024 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_95
timestamp 1679581782
transform 1 0 9696 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_102
timestamp 1679581782
transform 1 0 10368 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_109
timestamp 1679581782
transform 1 0 11040 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_116
timestamp 1679581782
transform 1 0 11712 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_123
timestamp 1679581782
transform 1 0 12384 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_130
timestamp 1679581782
transform 1 0 13056 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_137
timestamp 1679581782
transform 1 0 13728 0 1 21924
box -48 -56 720 834
use sg13g2_decap_4  FILLER_28_144
timestamp 1679577901
transform 1 0 14400 0 1 21924
box -48 -56 432 834
use sg13g2_fill_1  FILLER_28_148
timestamp 1677579658
transform 1 0 14784 0 1 21924
box -48 -56 144 834
use sg13g2_decap_8  FILLER_28_176
timestamp 1679581782
transform 1 0 17472 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_183
timestamp 1679581782
transform 1 0 18144 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_190
timestamp 1679581782
transform 1 0 18816 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_197
timestamp 1679581782
transform 1 0 19488 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_204
timestamp 1679581782
transform 1 0 20160 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_211
timestamp 1679581782
transform 1 0 20832 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_218
timestamp 1679581782
transform 1 0 21504 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_225
timestamp 1679581782
transform 1 0 22176 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_232
timestamp 1679581782
transform 1 0 22848 0 1 21924
box -48 -56 720 834
use sg13g2_decap_4  FILLER_28_239
timestamp 1679577901
transform 1 0 23520 0 1 21924
box -48 -56 432 834
use sg13g2_fill_2  FILLER_28_243
timestamp 1677580104
transform 1 0 23904 0 1 21924
box -48 -56 240 834
use sg13g2_decap_8  FILLER_28_272
timestamp 1679581782
transform 1 0 26688 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_279
timestamp 1679581782
transform 1 0 27360 0 1 21924
box -48 -56 720 834
use sg13g2_decap_4  FILLER_28_286
timestamp 1679577901
transform 1 0 28032 0 1 21924
box -48 -56 432 834
use sg13g2_fill_2  FILLER_28_290
timestamp 1677580104
transform 1 0 28416 0 1 21924
box -48 -56 240 834
use sg13g2_decap_8  FILLER_28_300
timestamp 1679581782
transform 1 0 29376 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_307
timestamp 1679581782
transform 1 0 30048 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_314
timestamp 1679581782
transform 1 0 30720 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_321
timestamp 1679581782
transform 1 0 31392 0 1 21924
box -48 -56 720 834
use sg13g2_fill_2  FILLER_28_328
timestamp 1677580104
transform 1 0 32064 0 1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_28_330
timestamp 1677579658
transform 1 0 32256 0 1 21924
box -48 -56 144 834
use sg13g2_decap_8  FILLER_28_335
timestamp 1679581782
transform 1 0 32736 0 1 21924
box -48 -56 720 834
use sg13g2_decap_4  FILLER_28_342
timestamp 1679577901
transform 1 0 33408 0 1 21924
box -48 -56 432 834
use sg13g2_fill_2  FILLER_28_346
timestamp 1677580104
transform 1 0 33792 0 1 21924
box -48 -56 240 834
use sg13g2_decap_8  FILLER_28_368
timestamp 1679581782
transform 1 0 35904 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_375
timestamp 1679581782
transform 1 0 36576 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_382
timestamp 1679581782
transform 1 0 37248 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_389
timestamp 1679581782
transform 1 0 37920 0 1 21924
box -48 -56 720 834
use sg13g2_decap_4  FILLER_28_396
timestamp 1679577901
transform 1 0 38592 0 1 21924
box -48 -56 432 834
use sg13g2_fill_1  FILLER_28_400
timestamp 1677579658
transform 1 0 38976 0 1 21924
box -48 -56 144 834
use sg13g2_decap_8  FILLER_28_428
timestamp 1679581782
transform 1 0 41664 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_435
timestamp 1679581782
transform 1 0 42336 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_442
timestamp 1679581782
transform 1 0 43008 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_449
timestamp 1679581782
transform 1 0 43680 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_456
timestamp 1679581782
transform 1 0 44352 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_463
timestamp 1679581782
transform 1 0 45024 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_470
timestamp 1679581782
transform 1 0 45696 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_477
timestamp 1679581782
transform 1 0 46368 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_484
timestamp 1679581782
transform 1 0 47040 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_491
timestamp 1679581782
transform 1 0 47712 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_498
timestamp 1679581782
transform 1 0 48384 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_505
timestamp 1679581782
transform 1 0 49056 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_512
timestamp 1679581782
transform 1 0 49728 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_519
timestamp 1679581782
transform 1 0 50400 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_526
timestamp 1679581782
transform 1 0 51072 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_533
timestamp 1679581782
transform 1 0 51744 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_540
timestamp 1679581782
transform 1 0 52416 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_547
timestamp 1679581782
transform 1 0 53088 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_554
timestamp 1679581782
transform 1 0 53760 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_561
timestamp 1679581782
transform 1 0 54432 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_568
timestamp 1679581782
transform 1 0 55104 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_575
timestamp 1679581782
transform 1 0 55776 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_582
timestamp 1679581782
transform 1 0 56448 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_589
timestamp 1679581782
transform 1 0 57120 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_596
timestamp 1679581782
transform 1 0 57792 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_603
timestamp 1679581782
transform 1 0 58464 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_610
timestamp 1679581782
transform 1 0 59136 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_617
timestamp 1679581782
transform 1 0 59808 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_624
timestamp 1679581782
transform 1 0 60480 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_631
timestamp 1679581782
transform 1 0 61152 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_638
timestamp 1679581782
transform 1 0 61824 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_645
timestamp 1679581782
transform 1 0 62496 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_652
timestamp 1679581782
transform 1 0 63168 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_659
timestamp 1679581782
transform 1 0 63840 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_666
timestamp 1679581782
transform 1 0 64512 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_673
timestamp 1679581782
transform 1 0 65184 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_680
timestamp 1679581782
transform 1 0 65856 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_687
timestamp 1679581782
transform 1 0 66528 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_694
timestamp 1679581782
transform 1 0 67200 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_701
timestamp 1679581782
transform 1 0 67872 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_708
timestamp 1679581782
transform 1 0 68544 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_715
timestamp 1679581782
transform 1 0 69216 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_722
timestamp 1679581782
transform 1 0 69888 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_729
timestamp 1679581782
transform 1 0 70560 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_736
timestamp 1679581782
transform 1 0 71232 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_743
timestamp 1679581782
transform 1 0 71904 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_750
timestamp 1679581782
transform 1 0 72576 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_757
timestamp 1679581782
transform 1 0 73248 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_764
timestamp 1679581782
transform 1 0 73920 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_771
timestamp 1679581782
transform 1 0 74592 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_778
timestamp 1679581782
transform 1 0 75264 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_785
timestamp 1679581782
transform 1 0 75936 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_792
timestamp 1679581782
transform 1 0 76608 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_799
timestamp 1679581782
transform 1 0 77280 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_806
timestamp 1679581782
transform 1 0 77952 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_813
timestamp 1679581782
transform 1 0 78624 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_820
timestamp 1679581782
transform 1 0 79296 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_827
timestamp 1679581782
transform 1 0 79968 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_834
timestamp 1679581782
transform 1 0 80640 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_841
timestamp 1679581782
transform 1 0 81312 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_848
timestamp 1679581782
transform 1 0 81984 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_855
timestamp 1679581782
transform 1 0 82656 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_862
timestamp 1679581782
transform 1 0 83328 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_869
timestamp 1679581782
transform 1 0 84000 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_876
timestamp 1679581782
transform 1 0 84672 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_883
timestamp 1679581782
transform 1 0 85344 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_890
timestamp 1679581782
transform 1 0 86016 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_897
timestamp 1679581782
transform 1 0 86688 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_904
timestamp 1679581782
transform 1 0 87360 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_911
timestamp 1679581782
transform 1 0 88032 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_918
timestamp 1679581782
transform 1 0 88704 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_925
timestamp 1679581782
transform 1 0 89376 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_932
timestamp 1679581782
transform 1 0 90048 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_939
timestamp 1679581782
transform 1 0 90720 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_946
timestamp 1679581782
transform 1 0 91392 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_953
timestamp 1679581782
transform 1 0 92064 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_960
timestamp 1679581782
transform 1 0 92736 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_967
timestamp 1679581782
transform 1 0 93408 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_974
timestamp 1679581782
transform 1 0 94080 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_981
timestamp 1679581782
transform 1 0 94752 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_988
timestamp 1679581782
transform 1 0 95424 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_995
timestamp 1679581782
transform 1 0 96096 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_1002
timestamp 1679581782
transform 1 0 96768 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_1009
timestamp 1679581782
transform 1 0 97440 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_1016
timestamp 1679581782
transform 1 0 98112 0 1 21924
box -48 -56 720 834
use sg13g2_decap_4  FILLER_28_1023
timestamp 1679577901
transform 1 0 98784 0 1 21924
box -48 -56 432 834
use sg13g2_fill_2  FILLER_28_1027
timestamp 1677580104
transform 1 0 99168 0 1 21924
box -48 -56 240 834
use sg13g2_decap_8  FILLER_29_0
timestamp 1679581782
transform 1 0 576 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_7
timestamp 1679581782
transform 1 0 1248 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_14
timestamp 1679581782
transform 1 0 1920 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_21
timestamp 1679581782
transform 1 0 2592 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_28
timestamp 1679581782
transform 1 0 3264 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_35
timestamp 1679581782
transform 1 0 3936 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_42
timestamp 1679581782
transform 1 0 4608 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_49
timestamp 1679581782
transform 1 0 5280 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_56
timestamp 1679581782
transform 1 0 5952 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_63
timestamp 1679581782
transform 1 0 6624 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_70
timestamp 1679581782
transform 1 0 7296 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_77
timestamp 1679581782
transform 1 0 7968 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_84
timestamp 1679581782
transform 1 0 8640 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_91
timestamp 1679581782
transform 1 0 9312 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_98
timestamp 1679581782
transform 1 0 9984 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_105
timestamp 1679581782
transform 1 0 10656 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_112
timestamp 1679581782
transform 1 0 11328 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_119
timestamp 1679581782
transform 1 0 12000 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_126
timestamp 1679581782
transform 1 0 12672 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_133
timestamp 1679581782
transform 1 0 13344 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_140
timestamp 1679581782
transform 1 0 14016 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_147
timestamp 1679581782
transform 1 0 14688 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_154
timestamp 1679581782
transform 1 0 15360 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_161
timestamp 1679581782
transform 1 0 16032 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_168
timestamp 1679581782
transform 1 0 16704 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_175
timestamp 1679581782
transform 1 0 17376 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_182
timestamp 1679581782
transform 1 0 18048 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_4  FILLER_29_189
timestamp 1679577901
transform 1 0 18720 0 -1 23436
box -48 -56 432 834
use sg13g2_fill_2  FILLER_29_193
timestamp 1677580104
transform 1 0 19104 0 -1 23436
box -48 -56 240 834
use sg13g2_decap_8  FILLER_29_222
timestamp 1679581782
transform 1 0 21888 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_229
timestamp 1679581782
transform 1 0 22560 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_236
timestamp 1679581782
transform 1 0 23232 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_243
timestamp 1679581782
transform 1 0 23904 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_250
timestamp 1679581782
transform 1 0 24576 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_257
timestamp 1679581782
transform 1 0 25248 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_264
timestamp 1679581782
transform 1 0 25920 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_271
timestamp 1679581782
transform 1 0 26592 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_278
timestamp 1679581782
transform 1 0 27264 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_4  FILLER_29_285
timestamp 1679577901
transform 1 0 27936 0 -1 23436
box -48 -56 432 834
use sg13g2_fill_2  FILLER_29_289
timestamp 1677580104
transform 1 0 28320 0 -1 23436
box -48 -56 240 834
use sg13g2_decap_8  FILLER_29_296
timestamp 1679581782
transform 1 0 28992 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_303
timestamp 1679581782
transform 1 0 29664 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_310
timestamp 1679581782
transform 1 0 30336 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_317
timestamp 1679581782
transform 1 0 31008 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_324
timestamp 1679581782
transform 1 0 31680 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_331
timestamp 1679581782
transform 1 0 32352 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_338
timestamp 1679581782
transform 1 0 33024 0 -1 23436
box -48 -56 720 834
use sg13g2_fill_2  FILLER_29_345
timestamp 1677580104
transform 1 0 33696 0 -1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_29_347
timestamp 1677579658
transform 1 0 33888 0 -1 23436
box -48 -56 144 834
use sg13g2_decap_8  FILLER_29_375
timestamp 1679581782
transform 1 0 36576 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_382
timestamp 1679581782
transform 1 0 37248 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_389
timestamp 1679581782
transform 1 0 37920 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_396
timestamp 1679581782
transform 1 0 38592 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_403
timestamp 1679581782
transform 1 0 39264 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_410
timestamp 1679581782
transform 1 0 39936 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_417
timestamp 1679581782
transform 1 0 40608 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_424
timestamp 1679581782
transform 1 0 41280 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_431
timestamp 1679581782
transform 1 0 41952 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_438
timestamp 1679581782
transform 1 0 42624 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_445
timestamp 1679581782
transform 1 0 43296 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_452
timestamp 1679581782
transform 1 0 43968 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_459
timestamp 1679581782
transform 1 0 44640 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_466
timestamp 1679581782
transform 1 0 45312 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_473
timestamp 1679581782
transform 1 0 45984 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_480
timestamp 1679581782
transform 1 0 46656 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_487
timestamp 1679581782
transform 1 0 47328 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_494
timestamp 1679581782
transform 1 0 48000 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_501
timestamp 1679581782
transform 1 0 48672 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_508
timestamp 1679581782
transform 1 0 49344 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_515
timestamp 1679581782
transform 1 0 50016 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_522
timestamp 1679581782
transform 1 0 50688 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_529
timestamp 1679581782
transform 1 0 51360 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_536
timestamp 1679581782
transform 1 0 52032 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_543
timestamp 1679581782
transform 1 0 52704 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_550
timestamp 1679581782
transform 1 0 53376 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_557
timestamp 1679581782
transform 1 0 54048 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_564
timestamp 1679581782
transform 1 0 54720 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_571
timestamp 1679581782
transform 1 0 55392 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_578
timestamp 1679581782
transform 1 0 56064 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_585
timestamp 1679581782
transform 1 0 56736 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_592
timestamp 1679581782
transform 1 0 57408 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_599
timestamp 1679581782
transform 1 0 58080 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_606
timestamp 1679581782
transform 1 0 58752 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_613
timestamp 1679581782
transform 1 0 59424 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_620
timestamp 1679581782
transform 1 0 60096 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_627
timestamp 1679581782
transform 1 0 60768 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_634
timestamp 1679581782
transform 1 0 61440 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_641
timestamp 1679581782
transform 1 0 62112 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_648
timestamp 1679581782
transform 1 0 62784 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_655
timestamp 1679581782
transform 1 0 63456 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_662
timestamp 1679581782
transform 1 0 64128 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_669
timestamp 1679581782
transform 1 0 64800 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_676
timestamp 1679581782
transform 1 0 65472 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_683
timestamp 1679581782
transform 1 0 66144 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_690
timestamp 1679581782
transform 1 0 66816 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_697
timestamp 1679581782
transform 1 0 67488 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_704
timestamp 1679581782
transform 1 0 68160 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_711
timestamp 1679581782
transform 1 0 68832 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_718
timestamp 1679581782
transform 1 0 69504 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_725
timestamp 1679581782
transform 1 0 70176 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_732
timestamp 1679581782
transform 1 0 70848 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_739
timestamp 1679581782
transform 1 0 71520 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_746
timestamp 1679581782
transform 1 0 72192 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_753
timestamp 1679581782
transform 1 0 72864 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_760
timestamp 1679581782
transform 1 0 73536 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_767
timestamp 1679581782
transform 1 0 74208 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_774
timestamp 1679581782
transform 1 0 74880 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_781
timestamp 1679581782
transform 1 0 75552 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_788
timestamp 1679581782
transform 1 0 76224 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_795
timestamp 1679581782
transform 1 0 76896 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_802
timestamp 1679581782
transform 1 0 77568 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_809
timestamp 1679581782
transform 1 0 78240 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_816
timestamp 1679581782
transform 1 0 78912 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_823
timestamp 1679581782
transform 1 0 79584 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_830
timestamp 1679581782
transform 1 0 80256 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_837
timestamp 1679581782
transform 1 0 80928 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_844
timestamp 1679581782
transform 1 0 81600 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_851
timestamp 1679581782
transform 1 0 82272 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_858
timestamp 1679581782
transform 1 0 82944 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_865
timestamp 1679581782
transform 1 0 83616 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_872
timestamp 1679581782
transform 1 0 84288 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_879
timestamp 1679581782
transform 1 0 84960 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_886
timestamp 1679581782
transform 1 0 85632 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_893
timestamp 1679581782
transform 1 0 86304 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_900
timestamp 1679581782
transform 1 0 86976 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_907
timestamp 1679581782
transform 1 0 87648 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_914
timestamp 1679581782
transform 1 0 88320 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_921
timestamp 1679581782
transform 1 0 88992 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_928
timestamp 1679581782
transform 1 0 89664 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_935
timestamp 1679581782
transform 1 0 90336 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_942
timestamp 1679581782
transform 1 0 91008 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_949
timestamp 1679581782
transform 1 0 91680 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_956
timestamp 1679581782
transform 1 0 92352 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_963
timestamp 1679581782
transform 1 0 93024 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_970
timestamp 1679581782
transform 1 0 93696 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_977
timestamp 1679581782
transform 1 0 94368 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_984
timestamp 1679581782
transform 1 0 95040 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_991
timestamp 1679581782
transform 1 0 95712 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_998
timestamp 1679581782
transform 1 0 96384 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_1005
timestamp 1679581782
transform 1 0 97056 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_1012
timestamp 1679581782
transform 1 0 97728 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_1019
timestamp 1679581782
transform 1 0 98400 0 -1 23436
box -48 -56 720 834
use sg13g2_fill_2  FILLER_29_1026
timestamp 1677580104
transform 1 0 99072 0 -1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_29_1028
timestamp 1677579658
transform 1 0 99264 0 -1 23436
box -48 -56 144 834
use sg13g2_decap_8  FILLER_30_5
timestamp 1679581782
transform 1 0 1056 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_12
timestamp 1679581782
transform 1 0 1728 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_19
timestamp 1679581782
transform 1 0 2400 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_26
timestamp 1679581782
transform 1 0 3072 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_33
timestamp 1679581782
transform 1 0 3744 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_40
timestamp 1679581782
transform 1 0 4416 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_47
timestamp 1679581782
transform 1 0 5088 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_54
timestamp 1679581782
transform 1 0 5760 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_61
timestamp 1679581782
transform 1 0 6432 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_68
timestamp 1679581782
transform 1 0 7104 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_75
timestamp 1679581782
transform 1 0 7776 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_82
timestamp 1679581782
transform 1 0 8448 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_89
timestamp 1679581782
transform 1 0 9120 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_96
timestamp 1679581782
transform 1 0 9792 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_103
timestamp 1679581782
transform 1 0 10464 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_110
timestamp 1679581782
transform 1 0 11136 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_117
timestamp 1679581782
transform 1 0 11808 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_124
timestamp 1679581782
transform 1 0 12480 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_131
timestamp 1679581782
transform 1 0 13152 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_138
timestamp 1679581782
transform 1 0 13824 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_145
timestamp 1679581782
transform 1 0 14496 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_152
timestamp 1679581782
transform 1 0 15168 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_159
timestamp 1679581782
transform 1 0 15840 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_166
timestamp 1679581782
transform 1 0 16512 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_173
timestamp 1679581782
transform 1 0 17184 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_180
timestamp 1679581782
transform 1 0 17856 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_187
timestamp 1679581782
transform 1 0 18528 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_194
timestamp 1679581782
transform 1 0 19200 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_201
timestamp 1679581782
transform 1 0 19872 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_208
timestamp 1679581782
transform 1 0 20544 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_215
timestamp 1679581782
transform 1 0 21216 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_222
timestamp 1679581782
transform 1 0 21888 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_229
timestamp 1679581782
transform 1 0 22560 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_236
timestamp 1679581782
transform 1 0 23232 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_243
timestamp 1679581782
transform 1 0 23904 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_250
timestamp 1679581782
transform 1 0 24576 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_257
timestamp 1679581782
transform 1 0 25248 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_264
timestamp 1679581782
transform 1 0 25920 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_271
timestamp 1679581782
transform 1 0 26592 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_278
timestamp 1679581782
transform 1 0 27264 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_285
timestamp 1679581782
transform 1 0 27936 0 1 23436
box -48 -56 720 834
use sg13g2_fill_2  FILLER_30_292
timestamp 1677580104
transform 1 0 28608 0 1 23436
box -48 -56 240 834
use sg13g2_decap_8  FILLER_30_297
timestamp 1679581782
transform 1 0 29088 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_304
timestamp 1679581782
transform 1 0 29760 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_311
timestamp 1679581782
transform 1 0 30432 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_318
timestamp 1679581782
transform 1 0 31104 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_325
timestamp 1679581782
transform 1 0 31776 0 1 23436
box -48 -56 720 834
use sg13g2_fill_2  FILLER_30_332
timestamp 1677580104
transform 1 0 32448 0 1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_30_334
timestamp 1677579658
transform 1 0 32640 0 1 23436
box -48 -56 144 834
use sg13g2_decap_8  FILLER_30_352
timestamp 1679581782
transform 1 0 34368 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_359
timestamp 1679581782
transform 1 0 35040 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_366
timestamp 1679581782
transform 1 0 35712 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_373
timestamp 1679581782
transform 1 0 36384 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_380
timestamp 1679581782
transform 1 0 37056 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_387
timestamp 1679581782
transform 1 0 37728 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_394
timestamp 1679581782
transform 1 0 38400 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_401
timestamp 1679581782
transform 1 0 39072 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_408
timestamp 1679581782
transform 1 0 39744 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_415
timestamp 1679581782
transform 1 0 40416 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_422
timestamp 1679581782
transform 1 0 41088 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_429
timestamp 1679581782
transform 1 0 41760 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_436
timestamp 1679581782
transform 1 0 42432 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_443
timestamp 1679581782
transform 1 0 43104 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_450
timestamp 1679581782
transform 1 0 43776 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_457
timestamp 1679581782
transform 1 0 44448 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_464
timestamp 1679581782
transform 1 0 45120 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_471
timestamp 1679581782
transform 1 0 45792 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_478
timestamp 1679581782
transform 1 0 46464 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_485
timestamp 1679581782
transform 1 0 47136 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_492
timestamp 1679581782
transform 1 0 47808 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_499
timestamp 1679581782
transform 1 0 48480 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_506
timestamp 1679581782
transform 1 0 49152 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_513
timestamp 1679581782
transform 1 0 49824 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_520
timestamp 1679581782
transform 1 0 50496 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_527
timestamp 1679581782
transform 1 0 51168 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_534
timestamp 1679581782
transform 1 0 51840 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_541
timestamp 1679581782
transform 1 0 52512 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_548
timestamp 1679581782
transform 1 0 53184 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_555
timestamp 1679581782
transform 1 0 53856 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_562
timestamp 1679581782
transform 1 0 54528 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_569
timestamp 1679581782
transform 1 0 55200 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_576
timestamp 1679581782
transform 1 0 55872 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_583
timestamp 1679581782
transform 1 0 56544 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_590
timestamp 1679581782
transform 1 0 57216 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_597
timestamp 1679581782
transform 1 0 57888 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_604
timestamp 1679581782
transform 1 0 58560 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_611
timestamp 1679581782
transform 1 0 59232 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_618
timestamp 1679581782
transform 1 0 59904 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_625
timestamp 1679581782
transform 1 0 60576 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_632
timestamp 1679581782
transform 1 0 61248 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_639
timestamp 1679581782
transform 1 0 61920 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_646
timestamp 1679581782
transform 1 0 62592 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_653
timestamp 1679581782
transform 1 0 63264 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_660
timestamp 1679581782
transform 1 0 63936 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_667
timestamp 1679581782
transform 1 0 64608 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_674
timestamp 1679581782
transform 1 0 65280 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_681
timestamp 1679581782
transform 1 0 65952 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_688
timestamp 1679581782
transform 1 0 66624 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_695
timestamp 1679581782
transform 1 0 67296 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_702
timestamp 1679581782
transform 1 0 67968 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_709
timestamp 1679581782
transform 1 0 68640 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_716
timestamp 1679581782
transform 1 0 69312 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_723
timestamp 1679581782
transform 1 0 69984 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_730
timestamp 1679581782
transform 1 0 70656 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_737
timestamp 1679581782
transform 1 0 71328 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_744
timestamp 1679581782
transform 1 0 72000 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_751
timestamp 1679581782
transform 1 0 72672 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_758
timestamp 1679581782
transform 1 0 73344 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_765
timestamp 1679581782
transform 1 0 74016 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_772
timestamp 1679581782
transform 1 0 74688 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_779
timestamp 1679581782
transform 1 0 75360 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_786
timestamp 1679581782
transform 1 0 76032 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_793
timestamp 1679581782
transform 1 0 76704 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_800
timestamp 1679581782
transform 1 0 77376 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_807
timestamp 1679581782
transform 1 0 78048 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_814
timestamp 1679581782
transform 1 0 78720 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_821
timestamp 1679581782
transform 1 0 79392 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_828
timestamp 1679581782
transform 1 0 80064 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_835
timestamp 1679581782
transform 1 0 80736 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_842
timestamp 1679581782
transform 1 0 81408 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_849
timestamp 1679581782
transform 1 0 82080 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_856
timestamp 1679581782
transform 1 0 82752 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_863
timestamp 1679581782
transform 1 0 83424 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_870
timestamp 1679581782
transform 1 0 84096 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_877
timestamp 1679581782
transform 1 0 84768 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_884
timestamp 1679581782
transform 1 0 85440 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_891
timestamp 1679581782
transform 1 0 86112 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_898
timestamp 1679581782
transform 1 0 86784 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_905
timestamp 1679581782
transform 1 0 87456 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_912
timestamp 1679581782
transform 1 0 88128 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_919
timestamp 1679581782
transform 1 0 88800 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_926
timestamp 1679581782
transform 1 0 89472 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_933
timestamp 1679581782
transform 1 0 90144 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_940
timestamp 1679581782
transform 1 0 90816 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_947
timestamp 1679581782
transform 1 0 91488 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_954
timestamp 1679581782
transform 1 0 92160 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_961
timestamp 1679581782
transform 1 0 92832 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_968
timestamp 1679581782
transform 1 0 93504 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_975
timestamp 1679581782
transform 1 0 94176 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_982
timestamp 1679581782
transform 1 0 94848 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_989
timestamp 1679581782
transform 1 0 95520 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_996
timestamp 1679581782
transform 1 0 96192 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_1003
timestamp 1679581782
transform 1 0 96864 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_1010
timestamp 1679581782
transform 1 0 97536 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_1017
timestamp 1679581782
transform 1 0 98208 0 1 23436
box -48 -56 720 834
use sg13g2_decap_4  FILLER_30_1024
timestamp 1679577901
transform 1 0 98880 0 1 23436
box -48 -56 432 834
use sg13g2_fill_1  FILLER_30_1028
timestamp 1677579658
transform 1 0 99264 0 1 23436
box -48 -56 144 834
use sg13g2_decap_8  FILLER_31_5
timestamp 1679581782
transform 1 0 1056 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_12
timestamp 1679581782
transform 1 0 1728 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_19
timestamp 1679581782
transform 1 0 2400 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_26
timestamp 1679581782
transform 1 0 3072 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_33
timestamp 1679581782
transform 1 0 3744 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_40
timestamp 1679581782
transform 1 0 4416 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_47
timestamp 1679581782
transform 1 0 5088 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_54
timestamp 1679581782
transform 1 0 5760 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_61
timestamp 1679581782
transform 1 0 6432 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_68
timestamp 1679581782
transform 1 0 7104 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_75
timestamp 1679581782
transform 1 0 7776 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_82
timestamp 1679581782
transform 1 0 8448 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_89
timestamp 1679581782
transform 1 0 9120 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_96
timestamp 1679581782
transform 1 0 9792 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_103
timestamp 1679581782
transform 1 0 10464 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_110
timestamp 1679581782
transform 1 0 11136 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_117
timestamp 1679581782
transform 1 0 11808 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_124
timestamp 1679581782
transform 1 0 12480 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_131
timestamp 1679581782
transform 1 0 13152 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_138
timestamp 1679581782
transform 1 0 13824 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_145
timestamp 1679581782
transform 1 0 14496 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_152
timestamp 1679581782
transform 1 0 15168 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_159
timestamp 1679581782
transform 1 0 15840 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_166
timestamp 1679581782
transform 1 0 16512 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_173
timestamp 1679581782
transform 1 0 17184 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_180
timestamp 1679581782
transform 1 0 17856 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_187
timestamp 1679581782
transform 1 0 18528 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_194
timestamp 1679581782
transform 1 0 19200 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_201
timestamp 1679581782
transform 1 0 19872 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_208
timestamp 1679581782
transform 1 0 20544 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_215
timestamp 1679581782
transform 1 0 21216 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_222
timestamp 1679581782
transform 1 0 21888 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_246
timestamp 1679581782
transform 1 0 24192 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_253
timestamp 1679581782
transform 1 0 24864 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_260
timestamp 1679581782
transform 1 0 25536 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_267
timestamp 1679581782
transform 1 0 26208 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_274
timestamp 1679581782
transform 1 0 26880 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_281
timestamp 1679581782
transform 1 0 27552 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_288
timestamp 1679581782
transform 1 0 28224 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_295
timestamp 1679581782
transform 1 0 28896 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_309
timestamp 1679581782
transform 1 0 30240 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_316
timestamp 1679581782
transform 1 0 30912 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_323
timestamp 1679581782
transform 1 0 31584 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_330
timestamp 1679581782
transform 1 0 32256 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_337
timestamp 1679581782
transform 1 0 32928 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_344
timestamp 1679581782
transform 1 0 33600 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_351
timestamp 1679581782
transform 1 0 34272 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_358
timestamp 1679581782
transform 1 0 34944 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_365
timestamp 1679581782
transform 1 0 35616 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_372
timestamp 1679581782
transform 1 0 36288 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_379
timestamp 1679581782
transform 1 0 36960 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_386
timestamp 1679581782
transform 1 0 37632 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_393
timestamp 1679581782
transform 1 0 38304 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_400
timestamp 1679581782
transform 1 0 38976 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_407
timestamp 1679581782
transform 1 0 39648 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_414
timestamp 1679581782
transform 1 0 40320 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_421
timestamp 1679581782
transform 1 0 40992 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_428
timestamp 1679581782
transform 1 0 41664 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_435
timestamp 1679581782
transform 1 0 42336 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_442
timestamp 1679581782
transform 1 0 43008 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_449
timestamp 1679581782
transform 1 0 43680 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_456
timestamp 1679581782
transform 1 0 44352 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_463
timestamp 1679581782
transform 1 0 45024 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_470
timestamp 1679581782
transform 1 0 45696 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_477
timestamp 1679581782
transform 1 0 46368 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_484
timestamp 1679581782
transform 1 0 47040 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_491
timestamp 1679581782
transform 1 0 47712 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_498
timestamp 1679581782
transform 1 0 48384 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_505
timestamp 1679581782
transform 1 0 49056 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_512
timestamp 1679581782
transform 1 0 49728 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_519
timestamp 1679581782
transform 1 0 50400 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_526
timestamp 1679581782
transform 1 0 51072 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_533
timestamp 1679581782
transform 1 0 51744 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_540
timestamp 1679581782
transform 1 0 52416 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_547
timestamp 1679581782
transform 1 0 53088 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_554
timestamp 1679581782
transform 1 0 53760 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_561
timestamp 1679581782
transform 1 0 54432 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_568
timestamp 1679581782
transform 1 0 55104 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_575
timestamp 1679581782
transform 1 0 55776 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_582
timestamp 1679581782
transform 1 0 56448 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_589
timestamp 1679581782
transform 1 0 57120 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_596
timestamp 1679581782
transform 1 0 57792 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_603
timestamp 1679581782
transform 1 0 58464 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_610
timestamp 1679581782
transform 1 0 59136 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_617
timestamp 1679581782
transform 1 0 59808 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_624
timestamp 1679581782
transform 1 0 60480 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_631
timestamp 1679581782
transform 1 0 61152 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_638
timestamp 1679581782
transform 1 0 61824 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_645
timestamp 1679581782
transform 1 0 62496 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_652
timestamp 1679581782
transform 1 0 63168 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_659
timestamp 1679581782
transform 1 0 63840 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_666
timestamp 1679581782
transform 1 0 64512 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_673
timestamp 1679581782
transform 1 0 65184 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_680
timestamp 1679581782
transform 1 0 65856 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_687
timestamp 1679581782
transform 1 0 66528 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_694
timestamp 1679581782
transform 1 0 67200 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_701
timestamp 1679581782
transform 1 0 67872 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_708
timestamp 1679581782
transform 1 0 68544 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_715
timestamp 1679581782
transform 1 0 69216 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_722
timestamp 1679581782
transform 1 0 69888 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_729
timestamp 1679581782
transform 1 0 70560 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_736
timestamp 1679581782
transform 1 0 71232 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_743
timestamp 1679581782
transform 1 0 71904 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_750
timestamp 1679581782
transform 1 0 72576 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_757
timestamp 1679581782
transform 1 0 73248 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_764
timestamp 1679581782
transform 1 0 73920 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_771
timestamp 1679581782
transform 1 0 74592 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_778
timestamp 1679581782
transform 1 0 75264 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_785
timestamp 1679581782
transform 1 0 75936 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_792
timestamp 1679581782
transform 1 0 76608 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_799
timestamp 1679581782
transform 1 0 77280 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_806
timestamp 1679581782
transform 1 0 77952 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_813
timestamp 1679581782
transform 1 0 78624 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_820
timestamp 1679581782
transform 1 0 79296 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_827
timestamp 1679581782
transform 1 0 79968 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_834
timestamp 1679581782
transform 1 0 80640 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_841
timestamp 1679581782
transform 1 0 81312 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_848
timestamp 1679581782
transform 1 0 81984 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_855
timestamp 1679581782
transform 1 0 82656 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_862
timestamp 1679581782
transform 1 0 83328 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_869
timestamp 1679581782
transform 1 0 84000 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_876
timestamp 1679581782
transform 1 0 84672 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_883
timestamp 1679581782
transform 1 0 85344 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_890
timestamp 1679581782
transform 1 0 86016 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_897
timestamp 1679581782
transform 1 0 86688 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_904
timestamp 1679581782
transform 1 0 87360 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_911
timestamp 1679581782
transform 1 0 88032 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_918
timestamp 1679581782
transform 1 0 88704 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_925
timestamp 1679581782
transform 1 0 89376 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_932
timestamp 1679581782
transform 1 0 90048 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_939
timestamp 1679581782
transform 1 0 90720 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_946
timestamp 1679581782
transform 1 0 91392 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_953
timestamp 1679581782
transform 1 0 92064 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_960
timestamp 1679581782
transform 1 0 92736 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_967
timestamp 1679581782
transform 1 0 93408 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_974
timestamp 1679581782
transform 1 0 94080 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_981
timestamp 1679581782
transform 1 0 94752 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_988
timestamp 1679581782
transform 1 0 95424 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_995
timestamp 1679581782
transform 1 0 96096 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_1002
timestamp 1679581782
transform 1 0 96768 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_1009
timestamp 1679581782
transform 1 0 97440 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_1016
timestamp 1679581782
transform 1 0 98112 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_4  FILLER_31_1023
timestamp 1679577901
transform 1 0 98784 0 -1 24948
box -48 -56 432 834
use sg13g2_fill_2  FILLER_31_1027
timestamp 1677580104
transform 1 0 99168 0 -1 24948
box -48 -56 240 834
use sg13g2_decap_8  FILLER_32_5
timestamp 1679581782
transform 1 0 1056 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_12
timestamp 1679581782
transform 1 0 1728 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_19
timestamp 1679581782
transform 1 0 2400 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_26
timestamp 1679581782
transform 1 0 3072 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_33
timestamp 1679581782
transform 1 0 3744 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_40
timestamp 1679581782
transform 1 0 4416 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_47
timestamp 1679581782
transform 1 0 5088 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_54
timestamp 1679581782
transform 1 0 5760 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_61
timestamp 1679581782
transform 1 0 6432 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_68
timestamp 1679581782
transform 1 0 7104 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_75
timestamp 1679581782
transform 1 0 7776 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_82
timestamp 1679581782
transform 1 0 8448 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_89
timestamp 1679581782
transform 1 0 9120 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_96
timestamp 1679581782
transform 1 0 9792 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_103
timestamp 1679581782
transform 1 0 10464 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_110
timestamp 1679581782
transform 1 0 11136 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_117
timestamp 1679581782
transform 1 0 11808 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_124
timestamp 1679581782
transform 1 0 12480 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_131
timestamp 1679581782
transform 1 0 13152 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_138
timestamp 1679581782
transform 1 0 13824 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_145
timestamp 1679581782
transform 1 0 14496 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_152
timestamp 1679581782
transform 1 0 15168 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_159
timestamp 1679581782
transform 1 0 15840 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_166
timestamp 1679581782
transform 1 0 16512 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_173
timestamp 1679581782
transform 1 0 17184 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_180
timestamp 1679581782
transform 1 0 17856 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_187
timestamp 1679581782
transform 1 0 18528 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_194
timestamp 1679581782
transform 1 0 19200 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_201
timestamp 1679581782
transform 1 0 19872 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_208
timestamp 1679581782
transform 1 0 20544 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_215
timestamp 1679581782
transform 1 0 21216 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_222
timestamp 1679581782
transform 1 0 21888 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_229
timestamp 1679581782
transform 1 0 22560 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_236
timestamp 1679581782
transform 1 0 23232 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_243
timestamp 1679581782
transform 1 0 23904 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_250
timestamp 1679581782
transform 1 0 24576 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_257
timestamp 1679581782
transform 1 0 25248 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_264
timestamp 1679581782
transform 1 0 25920 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_271
timestamp 1679581782
transform 1 0 26592 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_278
timestamp 1679581782
transform 1 0 27264 0 1 24948
box -48 -56 720 834
use sg13g2_fill_2  FILLER_32_285
timestamp 1677580104
transform 1 0 27936 0 1 24948
box -48 -56 240 834
use sg13g2_decap_8  FILLER_32_292
timestamp 1679581782
transform 1 0 28608 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_299
timestamp 1679581782
transform 1 0 29280 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_306
timestamp 1679581782
transform 1 0 29952 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_313
timestamp 1679581782
transform 1 0 30624 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_320
timestamp 1679581782
transform 1 0 31296 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_327
timestamp 1679581782
transform 1 0 31968 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_334
timestamp 1679581782
transform 1 0 32640 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_341
timestamp 1679581782
transform 1 0 33312 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_348
timestamp 1679581782
transform 1 0 33984 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_355
timestamp 1679581782
transform 1 0 34656 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_362
timestamp 1679581782
transform 1 0 35328 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_369
timestamp 1679581782
transform 1 0 36000 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_376
timestamp 1679581782
transform 1 0 36672 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_383
timestamp 1679581782
transform 1 0 37344 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_390
timestamp 1679581782
transform 1 0 38016 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_397
timestamp 1679581782
transform 1 0 38688 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_404
timestamp 1679581782
transform 1 0 39360 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_411
timestamp 1679581782
transform 1 0 40032 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_418
timestamp 1679581782
transform 1 0 40704 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_425
timestamp 1679581782
transform 1 0 41376 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_432
timestamp 1679581782
transform 1 0 42048 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_439
timestamp 1679581782
transform 1 0 42720 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_446
timestamp 1679581782
transform 1 0 43392 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_453
timestamp 1679581782
transform 1 0 44064 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_460
timestamp 1679581782
transform 1 0 44736 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_467
timestamp 1679581782
transform 1 0 45408 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_474
timestamp 1679581782
transform 1 0 46080 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_481
timestamp 1679581782
transform 1 0 46752 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_488
timestamp 1679581782
transform 1 0 47424 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_495
timestamp 1679581782
transform 1 0 48096 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_502
timestamp 1679581782
transform 1 0 48768 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_509
timestamp 1679581782
transform 1 0 49440 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_516
timestamp 1679581782
transform 1 0 50112 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_523
timestamp 1679581782
transform 1 0 50784 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_530
timestamp 1679581782
transform 1 0 51456 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_537
timestamp 1679581782
transform 1 0 52128 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_544
timestamp 1679581782
transform 1 0 52800 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_551
timestamp 1679581782
transform 1 0 53472 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_558
timestamp 1679581782
transform 1 0 54144 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_565
timestamp 1679581782
transform 1 0 54816 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_572
timestamp 1679581782
transform 1 0 55488 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_579
timestamp 1679581782
transform 1 0 56160 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_586
timestamp 1679581782
transform 1 0 56832 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_593
timestamp 1679581782
transform 1 0 57504 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_600
timestamp 1679581782
transform 1 0 58176 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_607
timestamp 1679581782
transform 1 0 58848 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_614
timestamp 1679581782
transform 1 0 59520 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_621
timestamp 1679581782
transform 1 0 60192 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_628
timestamp 1679581782
transform 1 0 60864 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_635
timestamp 1679581782
transform 1 0 61536 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_642
timestamp 1679581782
transform 1 0 62208 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_649
timestamp 1679581782
transform 1 0 62880 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_656
timestamp 1679581782
transform 1 0 63552 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_663
timestamp 1679581782
transform 1 0 64224 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_670
timestamp 1679581782
transform 1 0 64896 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_677
timestamp 1679581782
transform 1 0 65568 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_684
timestamp 1679581782
transform 1 0 66240 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_691
timestamp 1679581782
transform 1 0 66912 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_698
timestamp 1679581782
transform 1 0 67584 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_705
timestamp 1679581782
transform 1 0 68256 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_712
timestamp 1679581782
transform 1 0 68928 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_719
timestamp 1679581782
transform 1 0 69600 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_726
timestamp 1679581782
transform 1 0 70272 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_733
timestamp 1679581782
transform 1 0 70944 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_740
timestamp 1679581782
transform 1 0 71616 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_747
timestamp 1679581782
transform 1 0 72288 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_754
timestamp 1679581782
transform 1 0 72960 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_761
timestamp 1679581782
transform 1 0 73632 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_768
timestamp 1679581782
transform 1 0 74304 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_775
timestamp 1679581782
transform 1 0 74976 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_782
timestamp 1679581782
transform 1 0 75648 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_789
timestamp 1679581782
transform 1 0 76320 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_796
timestamp 1679581782
transform 1 0 76992 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_803
timestamp 1679581782
transform 1 0 77664 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_810
timestamp 1679581782
transform 1 0 78336 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_817
timestamp 1679581782
transform 1 0 79008 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_824
timestamp 1679581782
transform 1 0 79680 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_831
timestamp 1679581782
transform 1 0 80352 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_838
timestamp 1679581782
transform 1 0 81024 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_845
timestamp 1679581782
transform 1 0 81696 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_852
timestamp 1679581782
transform 1 0 82368 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_859
timestamp 1679581782
transform 1 0 83040 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_866
timestamp 1679581782
transform 1 0 83712 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_873
timestamp 1679581782
transform 1 0 84384 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_880
timestamp 1679581782
transform 1 0 85056 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_887
timestamp 1679581782
transform 1 0 85728 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_894
timestamp 1679581782
transform 1 0 86400 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_901
timestamp 1679581782
transform 1 0 87072 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_908
timestamp 1679581782
transform 1 0 87744 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_915
timestamp 1679581782
transform 1 0 88416 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_922
timestamp 1679581782
transform 1 0 89088 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_929
timestamp 1679581782
transform 1 0 89760 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_936
timestamp 1679581782
transform 1 0 90432 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_943
timestamp 1679581782
transform 1 0 91104 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_950
timestamp 1679581782
transform 1 0 91776 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_957
timestamp 1679581782
transform 1 0 92448 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_964
timestamp 1679581782
transform 1 0 93120 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_971
timestamp 1679581782
transform 1 0 93792 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_978
timestamp 1679581782
transform 1 0 94464 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_985
timestamp 1679581782
transform 1 0 95136 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_992
timestamp 1679581782
transform 1 0 95808 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_999
timestamp 1679581782
transform 1 0 96480 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_1006
timestamp 1679581782
transform 1 0 97152 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_1013
timestamp 1679581782
transform 1 0 97824 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_1020
timestamp 1679581782
transform 1 0 98496 0 1 24948
box -48 -56 720 834
use sg13g2_fill_2  FILLER_32_1027
timestamp 1677580104
transform 1 0 99168 0 1 24948
box -48 -56 240 834
use sg13g2_decap_8  FILLER_33_5
timestamp 1679581782
transform 1 0 1056 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_12
timestamp 1679581782
transform 1 0 1728 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_19
timestamp 1679581782
transform 1 0 2400 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_26
timestamp 1679581782
transform 1 0 3072 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_33
timestamp 1679581782
transform 1 0 3744 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_40
timestamp 1679581782
transform 1 0 4416 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_47
timestamp 1679581782
transform 1 0 5088 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_54
timestamp 1679581782
transform 1 0 5760 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_61
timestamp 1679581782
transform 1 0 6432 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_68
timestamp 1679581782
transform 1 0 7104 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_75
timestamp 1679581782
transform 1 0 7776 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_82
timestamp 1679581782
transform 1 0 8448 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_89
timestamp 1679581782
transform 1 0 9120 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_96
timestamp 1679581782
transform 1 0 9792 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_103
timestamp 1679581782
transform 1 0 10464 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_110
timestamp 1679581782
transform 1 0 11136 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_117
timestamp 1679581782
transform 1 0 11808 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_124
timestamp 1679581782
transform 1 0 12480 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_131
timestamp 1679581782
transform 1 0 13152 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_138
timestamp 1679581782
transform 1 0 13824 0 -1 26460
box -48 -56 720 834
use sg13g2_fill_2  FILLER_33_145
timestamp 1677580104
transform 1 0 14496 0 -1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_33_147
timestamp 1677579658
transform 1 0 14688 0 -1 26460
box -48 -56 144 834
use sg13g2_decap_8  FILLER_33_175
timestamp 1679581782
transform 1 0 17376 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_182
timestamp 1679581782
transform 1 0 18048 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_189
timestamp 1679581782
transform 1 0 18720 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_196
timestamp 1679581782
transform 1 0 19392 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_203
timestamp 1679581782
transform 1 0 20064 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_210
timestamp 1679581782
transform 1 0 20736 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_222
timestamp 1679581782
transform 1 0 21888 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_229
timestamp 1679581782
transform 1 0 22560 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_236
timestamp 1679581782
transform 1 0 23232 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_243
timestamp 1679581782
transform 1 0 23904 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_250
timestamp 1679581782
transform 1 0 24576 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_4  FILLER_33_257
timestamp 1679577901
transform 1 0 25248 0 -1 26460
box -48 -56 432 834
use sg13g2_fill_1  FILLER_33_261
timestamp 1677579658
transform 1 0 25632 0 -1 26460
box -48 -56 144 834
use sg13g2_decap_4  FILLER_33_279
timestamp 1679577901
transform 1 0 27360 0 -1 26460
box -48 -56 432 834
use sg13g2_fill_2  FILLER_33_283
timestamp 1677580104
transform 1 0 27744 0 -1 26460
box -48 -56 240 834
use sg13g2_decap_8  FILLER_33_291
timestamp 1679581782
transform 1 0 28512 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_298
timestamp 1679581782
transform 1 0 29184 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_305
timestamp 1679581782
transform 1 0 29856 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_312
timestamp 1679581782
transform 1 0 30528 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_319
timestamp 1679581782
transform 1 0 31200 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_326
timestamp 1679581782
transform 1 0 31872 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_333
timestamp 1679581782
transform 1 0 32544 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_340
timestamp 1679581782
transform 1 0 33216 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_4  FILLER_33_347
timestamp 1679577901
transform 1 0 33888 0 -1 26460
box -48 -56 432 834
use sg13g2_decap_8  FILLER_33_364
timestamp 1679581782
transform 1 0 35520 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_371
timestamp 1679581782
transform 1 0 36192 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_378
timestamp 1679581782
transform 1 0 36864 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_385
timestamp 1679581782
transform 1 0 37536 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_392
timestamp 1679581782
transform 1 0 38208 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_4  FILLER_33_399
timestamp 1679577901
transform 1 0 38880 0 -1 26460
box -48 -56 432 834
use sg13g2_fill_2  FILLER_33_403
timestamp 1677580104
transform 1 0 39264 0 -1 26460
box -48 -56 240 834
use sg13g2_decap_8  FILLER_33_418
timestamp 1679581782
transform 1 0 40704 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_425
timestamp 1679581782
transform 1 0 41376 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_432
timestamp 1679581782
transform 1 0 42048 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_439
timestamp 1679581782
transform 1 0 42720 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_446
timestamp 1679581782
transform 1 0 43392 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_453
timestamp 1679581782
transform 1 0 44064 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_460
timestamp 1679581782
transform 1 0 44736 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_467
timestamp 1679581782
transform 1 0 45408 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_474
timestamp 1679581782
transform 1 0 46080 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_481
timestamp 1679581782
transform 1 0 46752 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_488
timestamp 1679581782
transform 1 0 47424 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_495
timestamp 1679581782
transform 1 0 48096 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_502
timestamp 1679581782
transform 1 0 48768 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_509
timestamp 1679581782
transform 1 0 49440 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_516
timestamp 1679581782
transform 1 0 50112 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_523
timestamp 1679581782
transform 1 0 50784 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_530
timestamp 1679581782
transform 1 0 51456 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_537
timestamp 1679581782
transform 1 0 52128 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_544
timestamp 1679581782
transform 1 0 52800 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_551
timestamp 1679581782
transform 1 0 53472 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_558
timestamp 1679581782
transform 1 0 54144 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_565
timestamp 1679581782
transform 1 0 54816 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_572
timestamp 1679581782
transform 1 0 55488 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_579
timestamp 1679581782
transform 1 0 56160 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_586
timestamp 1679581782
transform 1 0 56832 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_593
timestamp 1679581782
transform 1 0 57504 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_600
timestamp 1679581782
transform 1 0 58176 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_607
timestamp 1679581782
transform 1 0 58848 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_614
timestamp 1679581782
transform 1 0 59520 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_621
timestamp 1679581782
transform 1 0 60192 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_628
timestamp 1679581782
transform 1 0 60864 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_635
timestamp 1679581782
transform 1 0 61536 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_642
timestamp 1679581782
transform 1 0 62208 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_649
timestamp 1679581782
transform 1 0 62880 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_656
timestamp 1679581782
transform 1 0 63552 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_663
timestamp 1679581782
transform 1 0 64224 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_670
timestamp 1679581782
transform 1 0 64896 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_677
timestamp 1679581782
transform 1 0 65568 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_684
timestamp 1679581782
transform 1 0 66240 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_691
timestamp 1679581782
transform 1 0 66912 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_698
timestamp 1679581782
transform 1 0 67584 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_705
timestamp 1679581782
transform 1 0 68256 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_712
timestamp 1679581782
transform 1 0 68928 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_719
timestamp 1679581782
transform 1 0 69600 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_726
timestamp 1679581782
transform 1 0 70272 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_733
timestamp 1679581782
transform 1 0 70944 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_740
timestamp 1679581782
transform 1 0 71616 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_747
timestamp 1679581782
transform 1 0 72288 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_754
timestamp 1679581782
transform 1 0 72960 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_761
timestamp 1679581782
transform 1 0 73632 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_768
timestamp 1679581782
transform 1 0 74304 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_775
timestamp 1679581782
transform 1 0 74976 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_782
timestamp 1679581782
transform 1 0 75648 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_789
timestamp 1679581782
transform 1 0 76320 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_796
timestamp 1679581782
transform 1 0 76992 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_803
timestamp 1679581782
transform 1 0 77664 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_810
timestamp 1679581782
transform 1 0 78336 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_817
timestamp 1679581782
transform 1 0 79008 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_824
timestamp 1679581782
transform 1 0 79680 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_831
timestamp 1679581782
transform 1 0 80352 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_838
timestamp 1679581782
transform 1 0 81024 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_845
timestamp 1679581782
transform 1 0 81696 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_852
timestamp 1679581782
transform 1 0 82368 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_859
timestamp 1679581782
transform 1 0 83040 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_866
timestamp 1679581782
transform 1 0 83712 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_873
timestamp 1679581782
transform 1 0 84384 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_880
timestamp 1679581782
transform 1 0 85056 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_887
timestamp 1679581782
transform 1 0 85728 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_894
timestamp 1679581782
transform 1 0 86400 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_901
timestamp 1679581782
transform 1 0 87072 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_908
timestamp 1679581782
transform 1 0 87744 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_915
timestamp 1679581782
transform 1 0 88416 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_922
timestamp 1679581782
transform 1 0 89088 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_929
timestamp 1679581782
transform 1 0 89760 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_936
timestamp 1679581782
transform 1 0 90432 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_943
timestamp 1679581782
transform 1 0 91104 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_950
timestamp 1679581782
transform 1 0 91776 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_957
timestamp 1679581782
transform 1 0 92448 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_964
timestamp 1679581782
transform 1 0 93120 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_971
timestamp 1679581782
transform 1 0 93792 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_978
timestamp 1679581782
transform 1 0 94464 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_985
timestamp 1679581782
transform 1 0 95136 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_992
timestamp 1679581782
transform 1 0 95808 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_999
timestamp 1679581782
transform 1 0 96480 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_1006
timestamp 1679581782
transform 1 0 97152 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_1013
timestamp 1679581782
transform 1 0 97824 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_1020
timestamp 1679581782
transform 1 0 98496 0 -1 26460
box -48 -56 720 834
use sg13g2_fill_2  FILLER_33_1027
timestamp 1677580104
transform 1 0 99168 0 -1 26460
box -48 -56 240 834
use sg13g2_decap_8  FILLER_34_5
timestamp 1679581782
transform 1 0 1056 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_12
timestamp 1679581782
transform 1 0 1728 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_19
timestamp 1679581782
transform 1 0 2400 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_26
timestamp 1679581782
transform 1 0 3072 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_33
timestamp 1679581782
transform 1 0 3744 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_40
timestamp 1679581782
transform 1 0 4416 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_47
timestamp 1679581782
transform 1 0 5088 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_54
timestamp 1679581782
transform 1 0 5760 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_61
timestamp 1679581782
transform 1 0 6432 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_68
timestamp 1679581782
transform 1 0 7104 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_75
timestamp 1679581782
transform 1 0 7776 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_82
timestamp 1679581782
transform 1 0 8448 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_89
timestamp 1679581782
transform 1 0 9120 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_96
timestamp 1679581782
transform 1 0 9792 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_103
timestamp 1679581782
transform 1 0 10464 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_110
timestamp 1679581782
transform 1 0 11136 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_117
timestamp 1679581782
transform 1 0 11808 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_124
timestamp 1679581782
transform 1 0 12480 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_131
timestamp 1679581782
transform 1 0 13152 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_138
timestamp 1679581782
transform 1 0 13824 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_145
timestamp 1679581782
transform 1 0 14496 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_152
timestamp 1679581782
transform 1 0 15168 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_159
timestamp 1679581782
transform 1 0 15840 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_166
timestamp 1679581782
transform 1 0 16512 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_173
timestamp 1679581782
transform 1 0 17184 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_180
timestamp 1679581782
transform 1 0 17856 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_187
timestamp 1679581782
transform 1 0 18528 0 1 26460
box -48 -56 720 834
use sg13g2_decap_4  FILLER_34_194
timestamp 1679577901
transform 1 0 19200 0 1 26460
box -48 -56 432 834
use sg13g2_fill_2  FILLER_34_198
timestamp 1677580104
transform 1 0 19584 0 1 26460
box -48 -56 240 834
use sg13g2_decap_8  FILLER_34_210
timestamp 1679581782
transform 1 0 20736 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_217
timestamp 1679581782
transform 1 0 21408 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_224
timestamp 1679581782
transform 1 0 22080 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_231
timestamp 1679581782
transform 1 0 22752 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_238
timestamp 1679581782
transform 1 0 23424 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_245
timestamp 1679581782
transform 1 0 24096 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_252
timestamp 1679581782
transform 1 0 24768 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_259
timestamp 1679581782
transform 1 0 25440 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_266
timestamp 1679581782
transform 1 0 26112 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_273
timestamp 1679581782
transform 1 0 26784 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_280
timestamp 1679581782
transform 1 0 27456 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_287
timestamp 1679581782
transform 1 0 28128 0 1 26460
box -48 -56 720 834
use sg13g2_decap_4  FILLER_34_294
timestamp 1679577901
transform 1 0 28800 0 1 26460
box -48 -56 432 834
use sg13g2_fill_2  FILLER_34_298
timestamp 1677580104
transform 1 0 29184 0 1 26460
box -48 -56 240 834
use sg13g2_decap_8  FILLER_34_310
timestamp 1679581782
transform 1 0 30336 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_317
timestamp 1679581782
transform 1 0 31008 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_324
timestamp 1679581782
transform 1 0 31680 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_331
timestamp 1679581782
transform 1 0 32352 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_338
timestamp 1679581782
transform 1 0 33024 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_345
timestamp 1679581782
transform 1 0 33696 0 1 26460
box -48 -56 720 834
use sg13g2_decap_4  FILLER_34_352
timestamp 1679577901
transform 1 0 34368 0 1 26460
box -48 -56 432 834
use sg13g2_fill_1  FILLER_34_356
timestamp 1677579658
transform 1 0 34752 0 1 26460
box -48 -56 144 834
use sg13g2_decap_8  FILLER_34_384
timestamp 1679581782
transform 1 0 37440 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_391
timestamp 1679581782
transform 1 0 38112 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_398
timestamp 1679581782
transform 1 0 38784 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_405
timestamp 1679581782
transform 1 0 39456 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_412
timestamp 1679581782
transform 1 0 40128 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_419
timestamp 1679581782
transform 1 0 40800 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_426
timestamp 1679581782
transform 1 0 41472 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_433
timestamp 1679581782
transform 1 0 42144 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_440
timestamp 1679581782
transform 1 0 42816 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_447
timestamp 1679581782
transform 1 0 43488 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_454
timestamp 1679581782
transform 1 0 44160 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_461
timestamp 1679581782
transform 1 0 44832 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_468
timestamp 1679581782
transform 1 0 45504 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_475
timestamp 1679581782
transform 1 0 46176 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_482
timestamp 1679581782
transform 1 0 46848 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_489
timestamp 1679581782
transform 1 0 47520 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_496
timestamp 1679581782
transform 1 0 48192 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_503
timestamp 1679581782
transform 1 0 48864 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_510
timestamp 1679581782
transform 1 0 49536 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_517
timestamp 1679581782
transform 1 0 50208 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_524
timestamp 1679581782
transform 1 0 50880 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_531
timestamp 1679581782
transform 1 0 51552 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_538
timestamp 1679581782
transform 1 0 52224 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_545
timestamp 1679581782
transform 1 0 52896 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_552
timestamp 1679581782
transform 1 0 53568 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_559
timestamp 1679581782
transform 1 0 54240 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_566
timestamp 1679581782
transform 1 0 54912 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_573
timestamp 1679581782
transform 1 0 55584 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_580
timestamp 1679581782
transform 1 0 56256 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_587
timestamp 1679581782
transform 1 0 56928 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_594
timestamp 1679581782
transform 1 0 57600 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_601
timestamp 1679581782
transform 1 0 58272 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_608
timestamp 1679581782
transform 1 0 58944 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_615
timestamp 1679581782
transform 1 0 59616 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_622
timestamp 1679581782
transform 1 0 60288 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_629
timestamp 1679581782
transform 1 0 60960 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_636
timestamp 1679581782
transform 1 0 61632 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_643
timestamp 1679581782
transform 1 0 62304 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_650
timestamp 1679581782
transform 1 0 62976 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_657
timestamp 1679581782
transform 1 0 63648 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_664
timestamp 1679581782
transform 1 0 64320 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_671
timestamp 1679581782
transform 1 0 64992 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_678
timestamp 1679581782
transform 1 0 65664 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_685
timestamp 1679581782
transform 1 0 66336 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_692
timestamp 1679581782
transform 1 0 67008 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_699
timestamp 1679581782
transform 1 0 67680 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_706
timestamp 1679581782
transform 1 0 68352 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_713
timestamp 1679581782
transform 1 0 69024 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_720
timestamp 1679581782
transform 1 0 69696 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_727
timestamp 1679581782
transform 1 0 70368 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_734
timestamp 1679581782
transform 1 0 71040 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_741
timestamp 1679581782
transform 1 0 71712 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_748
timestamp 1679581782
transform 1 0 72384 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_755
timestamp 1679581782
transform 1 0 73056 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_762
timestamp 1679581782
transform 1 0 73728 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_769
timestamp 1679581782
transform 1 0 74400 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_776
timestamp 1679581782
transform 1 0 75072 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_783
timestamp 1679581782
transform 1 0 75744 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_790
timestamp 1679581782
transform 1 0 76416 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_797
timestamp 1679581782
transform 1 0 77088 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_804
timestamp 1679581782
transform 1 0 77760 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_811
timestamp 1679581782
transform 1 0 78432 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_818
timestamp 1679581782
transform 1 0 79104 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_825
timestamp 1679581782
transform 1 0 79776 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_832
timestamp 1679581782
transform 1 0 80448 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_839
timestamp 1679581782
transform 1 0 81120 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_846
timestamp 1679581782
transform 1 0 81792 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_853
timestamp 1679581782
transform 1 0 82464 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_860
timestamp 1679581782
transform 1 0 83136 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_867
timestamp 1679581782
transform 1 0 83808 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_874
timestamp 1679581782
transform 1 0 84480 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_881
timestamp 1679581782
transform 1 0 85152 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_888
timestamp 1679581782
transform 1 0 85824 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_895
timestamp 1679581782
transform 1 0 86496 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_902
timestamp 1679581782
transform 1 0 87168 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_909
timestamp 1679581782
transform 1 0 87840 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_916
timestamp 1679581782
transform 1 0 88512 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_923
timestamp 1679581782
transform 1 0 89184 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_930
timestamp 1679581782
transform 1 0 89856 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_937
timestamp 1679581782
transform 1 0 90528 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_944
timestamp 1679581782
transform 1 0 91200 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_951
timestamp 1679581782
transform 1 0 91872 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_958
timestamp 1679581782
transform 1 0 92544 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_965
timestamp 1679581782
transform 1 0 93216 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_972
timestamp 1679581782
transform 1 0 93888 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_979
timestamp 1679581782
transform 1 0 94560 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_986
timestamp 1679581782
transform 1 0 95232 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_993
timestamp 1679581782
transform 1 0 95904 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_1000
timestamp 1679581782
transform 1 0 96576 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_1007
timestamp 1679581782
transform 1 0 97248 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_1014
timestamp 1679581782
transform 1 0 97920 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_1021
timestamp 1679581782
transform 1 0 98592 0 1 26460
box -48 -56 720 834
use sg13g2_fill_1  FILLER_34_1028
timestamp 1677579658
transform 1 0 99264 0 1 26460
box -48 -56 144 834
use sg13g2_decap_8  FILLER_35_5
timestamp 1679581782
transform 1 0 1056 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_12
timestamp 1679581782
transform 1 0 1728 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_19
timestamp 1679581782
transform 1 0 2400 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_26
timestamp 1679581782
transform 1 0 3072 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_33
timestamp 1679581782
transform 1 0 3744 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_40
timestamp 1679581782
transform 1 0 4416 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_47
timestamp 1679581782
transform 1 0 5088 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_54
timestamp 1679581782
transform 1 0 5760 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_61
timestamp 1679581782
transform 1 0 6432 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_68
timestamp 1679581782
transform 1 0 7104 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_75
timestamp 1679581782
transform 1 0 7776 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_82
timestamp 1679581782
transform 1 0 8448 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_89
timestamp 1679581782
transform 1 0 9120 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_96
timestamp 1679581782
transform 1 0 9792 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_103
timestamp 1679581782
transform 1 0 10464 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_110
timestamp 1679581782
transform 1 0 11136 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_117
timestamp 1679581782
transform 1 0 11808 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_124
timestamp 1679581782
transform 1 0 12480 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_131
timestamp 1679581782
transform 1 0 13152 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_138
timestamp 1679581782
transform 1 0 13824 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_145
timestamp 1679581782
transform 1 0 14496 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_152
timestamp 1679581782
transform 1 0 15168 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_159
timestamp 1679581782
transform 1 0 15840 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_166
timestamp 1679581782
transform 1 0 16512 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_173
timestamp 1679581782
transform 1 0 17184 0 -1 27972
box -48 -56 720 834
use sg13g2_fill_2  FILLER_35_180
timestamp 1677580104
transform 1 0 17856 0 -1 27972
box -48 -56 240 834
use sg13g2_decap_8  FILLER_35_192
timestamp 1679581782
transform 1 0 19008 0 -1 27972
box -48 -56 720 834
use sg13g2_fill_2  FILLER_35_199
timestamp 1677580104
transform 1 0 19680 0 -1 27972
box -48 -56 240 834
use sg13g2_fill_1  FILLER_35_201
timestamp 1677579658
transform 1 0 19872 0 -1 27972
box -48 -56 144 834
use sg13g2_decap_8  FILLER_35_207
timestamp 1679581782
transform 1 0 20448 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_214
timestamp 1679581782
transform 1 0 21120 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_221
timestamp 1679581782
transform 1 0 21792 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_228
timestamp 1679581782
transform 1 0 22464 0 -1 27972
box -48 -56 720 834
use sg13g2_fill_1  FILLER_35_235
timestamp 1677579658
transform 1 0 23136 0 -1 27972
box -48 -56 144 834
use sg13g2_decap_8  FILLER_35_241
timestamp 1679581782
transform 1 0 23712 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_248
timestamp 1679581782
transform 1 0 24384 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_255
timestamp 1679581782
transform 1 0 25056 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_4  FILLER_35_262
timestamp 1679577901
transform 1 0 25728 0 -1 27972
box -48 -56 432 834
use sg13g2_fill_2  FILLER_35_266
timestamp 1677580104
transform 1 0 26112 0 -1 27972
box -48 -56 240 834
use sg13g2_decap_8  FILLER_35_278
timestamp 1679581782
transform 1 0 27264 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_285
timestamp 1679581782
transform 1 0 27936 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_4  FILLER_35_292
timestamp 1679577901
transform 1 0 28608 0 -1 27972
box -48 -56 432 834
use sg13g2_fill_2  FILLER_35_296
timestamp 1677580104
transform 1 0 28992 0 -1 27972
box -48 -56 240 834
use sg13g2_decap_8  FILLER_35_304
timestamp 1679581782
transform 1 0 29760 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_311
timestamp 1679581782
transform 1 0 30432 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_318
timestamp 1679581782
transform 1 0 31104 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_325
timestamp 1679581782
transform 1 0 31776 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_332
timestamp 1679581782
transform 1 0 32448 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_339
timestamp 1679581782
transform 1 0 33120 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_346
timestamp 1679581782
transform 1 0 33792 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_353
timestamp 1679581782
transform 1 0 34464 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_360
timestamp 1679581782
transform 1 0 35136 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_367
timestamp 1679581782
transform 1 0 35808 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_374
timestamp 1679581782
transform 1 0 36480 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_381
timestamp 1679581782
transform 1 0 37152 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_388
timestamp 1679581782
transform 1 0 37824 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_395
timestamp 1679581782
transform 1 0 38496 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_402
timestamp 1679581782
transform 1 0 39168 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_409
timestamp 1679581782
transform 1 0 39840 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_416
timestamp 1679581782
transform 1 0 40512 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_423
timestamp 1679581782
transform 1 0 41184 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_430
timestamp 1679581782
transform 1 0 41856 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_437
timestamp 1679581782
transform 1 0 42528 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_444
timestamp 1679581782
transform 1 0 43200 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_451
timestamp 1679581782
transform 1 0 43872 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_458
timestamp 1679581782
transform 1 0 44544 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_465
timestamp 1679581782
transform 1 0 45216 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_472
timestamp 1679581782
transform 1 0 45888 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_479
timestamp 1679581782
transform 1 0 46560 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_486
timestamp 1679581782
transform 1 0 47232 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_493
timestamp 1679581782
transform 1 0 47904 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_500
timestamp 1679581782
transform 1 0 48576 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_507
timestamp 1679581782
transform 1 0 49248 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_514
timestamp 1679581782
transform 1 0 49920 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_521
timestamp 1679581782
transform 1 0 50592 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_528
timestamp 1679581782
transform 1 0 51264 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_535
timestamp 1679581782
transform 1 0 51936 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_542
timestamp 1679581782
transform 1 0 52608 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_549
timestamp 1679581782
transform 1 0 53280 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_556
timestamp 1679581782
transform 1 0 53952 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_563
timestamp 1679581782
transform 1 0 54624 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_570
timestamp 1679581782
transform 1 0 55296 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_577
timestamp 1679581782
transform 1 0 55968 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_584
timestamp 1679581782
transform 1 0 56640 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_591
timestamp 1679581782
transform 1 0 57312 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_598
timestamp 1679581782
transform 1 0 57984 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_605
timestamp 1679581782
transform 1 0 58656 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_612
timestamp 1679581782
transform 1 0 59328 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_619
timestamp 1679581782
transform 1 0 60000 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_626
timestamp 1679581782
transform 1 0 60672 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_633
timestamp 1679581782
transform 1 0 61344 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_640
timestamp 1679581782
transform 1 0 62016 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_647
timestamp 1679581782
transform 1 0 62688 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_654
timestamp 1679581782
transform 1 0 63360 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_661
timestamp 1679581782
transform 1 0 64032 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_668
timestamp 1679581782
transform 1 0 64704 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_675
timestamp 1679581782
transform 1 0 65376 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_682
timestamp 1679581782
transform 1 0 66048 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_689
timestamp 1679581782
transform 1 0 66720 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_696
timestamp 1679581782
transform 1 0 67392 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_703
timestamp 1679581782
transform 1 0 68064 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_710
timestamp 1679581782
transform 1 0 68736 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_717
timestamp 1679581782
transform 1 0 69408 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_724
timestamp 1679581782
transform 1 0 70080 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_731
timestamp 1679581782
transform 1 0 70752 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_738
timestamp 1679581782
transform 1 0 71424 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_745
timestamp 1679581782
transform 1 0 72096 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_752
timestamp 1679581782
transform 1 0 72768 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_759
timestamp 1679581782
transform 1 0 73440 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_766
timestamp 1679581782
transform 1 0 74112 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_773
timestamp 1679581782
transform 1 0 74784 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_780
timestamp 1679581782
transform 1 0 75456 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_787
timestamp 1679581782
transform 1 0 76128 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_794
timestamp 1679581782
transform 1 0 76800 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_801
timestamp 1679581782
transform 1 0 77472 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_808
timestamp 1679581782
transform 1 0 78144 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_815
timestamp 1679581782
transform 1 0 78816 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_822
timestamp 1679581782
transform 1 0 79488 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_829
timestamp 1679581782
transform 1 0 80160 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_836
timestamp 1679581782
transform 1 0 80832 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_843
timestamp 1679581782
transform 1 0 81504 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_850
timestamp 1679581782
transform 1 0 82176 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_857
timestamp 1679581782
transform 1 0 82848 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_864
timestamp 1679581782
transform 1 0 83520 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_871
timestamp 1679581782
transform 1 0 84192 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_878
timestamp 1679581782
transform 1 0 84864 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_885
timestamp 1679581782
transform 1 0 85536 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_892
timestamp 1679581782
transform 1 0 86208 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_899
timestamp 1679581782
transform 1 0 86880 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_906
timestamp 1679581782
transform 1 0 87552 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_913
timestamp 1679581782
transform 1 0 88224 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_920
timestamp 1679581782
transform 1 0 88896 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_927
timestamp 1679581782
transform 1 0 89568 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_934
timestamp 1679581782
transform 1 0 90240 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_941
timestamp 1679581782
transform 1 0 90912 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_948
timestamp 1679581782
transform 1 0 91584 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_955
timestamp 1679581782
transform 1 0 92256 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_962
timestamp 1679581782
transform 1 0 92928 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_969
timestamp 1679581782
transform 1 0 93600 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_976
timestamp 1679581782
transform 1 0 94272 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_983
timestamp 1679581782
transform 1 0 94944 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_990
timestamp 1679581782
transform 1 0 95616 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_997
timestamp 1679581782
transform 1 0 96288 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_1004
timestamp 1679581782
transform 1 0 96960 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_1011
timestamp 1679581782
transform 1 0 97632 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_1018
timestamp 1679581782
transform 1 0 98304 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_4  FILLER_35_1025
timestamp 1679577901
transform 1 0 98976 0 -1 27972
box -48 -56 432 834
use sg13g2_decap_8  FILLER_36_5
timestamp 1679581782
transform 1 0 1056 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_12
timestamp 1679581782
transform 1 0 1728 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_19
timestamp 1679581782
transform 1 0 2400 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_26
timestamp 1679581782
transform 1 0 3072 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_33
timestamp 1679581782
transform 1 0 3744 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_40
timestamp 1679581782
transform 1 0 4416 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_47
timestamp 1679581782
transform 1 0 5088 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_54
timestamp 1679581782
transform 1 0 5760 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_61
timestamp 1679581782
transform 1 0 6432 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_68
timestamp 1679581782
transform 1 0 7104 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_75
timestamp 1679581782
transform 1 0 7776 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_82
timestamp 1679581782
transform 1 0 8448 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_89
timestamp 1679581782
transform 1 0 9120 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_96
timestamp 1679581782
transform 1 0 9792 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_103
timestamp 1679581782
transform 1 0 10464 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_110
timestamp 1679581782
transform 1 0 11136 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_117
timestamp 1679581782
transform 1 0 11808 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_124
timestamp 1679581782
transform 1 0 12480 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_131
timestamp 1679581782
transform 1 0 13152 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_138
timestamp 1679581782
transform 1 0 13824 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_145
timestamp 1679581782
transform 1 0 14496 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_152
timestamp 1679581782
transform 1 0 15168 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_159
timestamp 1679581782
transform 1 0 15840 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_166
timestamp 1679581782
transform 1 0 16512 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_173
timestamp 1679581782
transform 1 0 17184 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_180
timestamp 1679581782
transform 1 0 17856 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_187
timestamp 1679581782
transform 1 0 18528 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_194
timestamp 1679581782
transform 1 0 19200 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_201
timestamp 1679581782
transform 1 0 19872 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_208
timestamp 1679581782
transform 1 0 20544 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_215
timestamp 1679581782
transform 1 0 21216 0 1 27972
box -48 -56 720 834
use sg13g2_fill_1  FILLER_36_222
timestamp 1677579658
transform 1 0 21888 0 1 27972
box -48 -56 144 834
use sg13g2_decap_4  FILLER_36_230
timestamp 1679577901
transform 1 0 22656 0 1 27972
box -48 -56 432 834
use sg13g2_fill_1  FILLER_36_234
timestamp 1677579658
transform 1 0 23040 0 1 27972
box -48 -56 144 834
use sg13g2_decap_8  FILLER_36_240
timestamp 1679581782
transform 1 0 23616 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_247
timestamp 1679581782
transform 1 0 24288 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_254
timestamp 1679581782
transform 1 0 24960 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_261
timestamp 1679581782
transform 1 0 25632 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_268
timestamp 1679581782
transform 1 0 26304 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_275
timestamp 1679581782
transform 1 0 26976 0 1 27972
box -48 -56 720 834
use sg13g2_decap_4  FILLER_36_282
timestamp 1679577901
transform 1 0 27648 0 1 27972
box -48 -56 432 834
use sg13g2_fill_1  FILLER_36_292
timestamp 1677579658
transform 1 0 28608 0 1 27972
box -48 -56 144 834
use sg13g2_decap_8  FILLER_36_305
timestamp 1679581782
transform 1 0 29856 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_312
timestamp 1679581782
transform 1 0 30528 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_319
timestamp 1679581782
transform 1 0 31200 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_326
timestamp 1679581782
transform 1 0 31872 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_333
timestamp 1679581782
transform 1 0 32544 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_340
timestamp 1679581782
transform 1 0 33216 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_347
timestamp 1679581782
transform 1 0 33888 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_354
timestamp 1679581782
transform 1 0 34560 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_361
timestamp 1679581782
transform 1 0 35232 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_368
timestamp 1679581782
transform 1 0 35904 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_375
timestamp 1679581782
transform 1 0 36576 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_382
timestamp 1679581782
transform 1 0 37248 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_389
timestamp 1679581782
transform 1 0 37920 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_396
timestamp 1679581782
transform 1 0 38592 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_403
timestamp 1679581782
transform 1 0 39264 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_410
timestamp 1679581782
transform 1 0 39936 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_417
timestamp 1679581782
transform 1 0 40608 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_424
timestamp 1679581782
transform 1 0 41280 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_431
timestamp 1679581782
transform 1 0 41952 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_438
timestamp 1679581782
transform 1 0 42624 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_445
timestamp 1679581782
transform 1 0 43296 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_452
timestamp 1679581782
transform 1 0 43968 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_459
timestamp 1679581782
transform 1 0 44640 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_466
timestamp 1679581782
transform 1 0 45312 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_473
timestamp 1679581782
transform 1 0 45984 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_480
timestamp 1679581782
transform 1 0 46656 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_487
timestamp 1679581782
transform 1 0 47328 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_494
timestamp 1679581782
transform 1 0 48000 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_501
timestamp 1679581782
transform 1 0 48672 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_508
timestamp 1679581782
transform 1 0 49344 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_515
timestamp 1679581782
transform 1 0 50016 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_522
timestamp 1679581782
transform 1 0 50688 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_529
timestamp 1679581782
transform 1 0 51360 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_536
timestamp 1679581782
transform 1 0 52032 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_543
timestamp 1679581782
transform 1 0 52704 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_550
timestamp 1679581782
transform 1 0 53376 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_557
timestamp 1679581782
transform 1 0 54048 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_564
timestamp 1679581782
transform 1 0 54720 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_571
timestamp 1679581782
transform 1 0 55392 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_578
timestamp 1679581782
transform 1 0 56064 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_585
timestamp 1679581782
transform 1 0 56736 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_592
timestamp 1679581782
transform 1 0 57408 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_599
timestamp 1679581782
transform 1 0 58080 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_606
timestamp 1679581782
transform 1 0 58752 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_613
timestamp 1679581782
transform 1 0 59424 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_620
timestamp 1679581782
transform 1 0 60096 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_627
timestamp 1679581782
transform 1 0 60768 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_634
timestamp 1679581782
transform 1 0 61440 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_641
timestamp 1679581782
transform 1 0 62112 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_648
timestamp 1679581782
transform 1 0 62784 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_655
timestamp 1679581782
transform 1 0 63456 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_662
timestamp 1679581782
transform 1 0 64128 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_669
timestamp 1679581782
transform 1 0 64800 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_676
timestamp 1679581782
transform 1 0 65472 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_683
timestamp 1679581782
transform 1 0 66144 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_690
timestamp 1679581782
transform 1 0 66816 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_697
timestamp 1679581782
transform 1 0 67488 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_704
timestamp 1679581782
transform 1 0 68160 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_711
timestamp 1679581782
transform 1 0 68832 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_718
timestamp 1679581782
transform 1 0 69504 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_725
timestamp 1679581782
transform 1 0 70176 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_732
timestamp 1679581782
transform 1 0 70848 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_739
timestamp 1679581782
transform 1 0 71520 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_746
timestamp 1679581782
transform 1 0 72192 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_753
timestamp 1679581782
transform 1 0 72864 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_760
timestamp 1679581782
transform 1 0 73536 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_767
timestamp 1679581782
transform 1 0 74208 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_774
timestamp 1679581782
transform 1 0 74880 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_781
timestamp 1679581782
transform 1 0 75552 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_788
timestamp 1679581782
transform 1 0 76224 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_795
timestamp 1679581782
transform 1 0 76896 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_802
timestamp 1679581782
transform 1 0 77568 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_809
timestamp 1679581782
transform 1 0 78240 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_816
timestamp 1679581782
transform 1 0 78912 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_823
timestamp 1679581782
transform 1 0 79584 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_830
timestamp 1679581782
transform 1 0 80256 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_837
timestamp 1679581782
transform 1 0 80928 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_844
timestamp 1679581782
transform 1 0 81600 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_851
timestamp 1679581782
transform 1 0 82272 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_858
timestamp 1679581782
transform 1 0 82944 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_865
timestamp 1679581782
transform 1 0 83616 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_872
timestamp 1679581782
transform 1 0 84288 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_879
timestamp 1679581782
transform 1 0 84960 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_886
timestamp 1679581782
transform 1 0 85632 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_893
timestamp 1679581782
transform 1 0 86304 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_900
timestamp 1679581782
transform 1 0 86976 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_907
timestamp 1679581782
transform 1 0 87648 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_914
timestamp 1679581782
transform 1 0 88320 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_921
timestamp 1679581782
transform 1 0 88992 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_928
timestamp 1679581782
transform 1 0 89664 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_935
timestamp 1679581782
transform 1 0 90336 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_942
timestamp 1679581782
transform 1 0 91008 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_949
timestamp 1679581782
transform 1 0 91680 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_956
timestamp 1679581782
transform 1 0 92352 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_963
timestamp 1679581782
transform 1 0 93024 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_970
timestamp 1679581782
transform 1 0 93696 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_977
timestamp 1679581782
transform 1 0 94368 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_984
timestamp 1679581782
transform 1 0 95040 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_991
timestamp 1679581782
transform 1 0 95712 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_998
timestamp 1679581782
transform 1 0 96384 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_1005
timestamp 1679581782
transform 1 0 97056 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_1012
timestamp 1679581782
transform 1 0 97728 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_1019
timestamp 1679581782
transform 1 0 98400 0 1 27972
box -48 -56 720 834
use sg13g2_fill_2  FILLER_36_1026
timestamp 1677580104
transform 1 0 99072 0 1 27972
box -48 -56 240 834
use sg13g2_fill_1  FILLER_36_1028
timestamp 1677579658
transform 1 0 99264 0 1 27972
box -48 -56 144 834
use sg13g2_decap_8  FILLER_37_0
timestamp 1679581782
transform 1 0 576 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_7
timestamp 1679581782
transform 1 0 1248 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_14
timestamp 1679581782
transform 1 0 1920 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_21
timestamp 1679581782
transform 1 0 2592 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_28
timestamp 1679581782
transform 1 0 3264 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_35
timestamp 1679581782
transform 1 0 3936 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_42
timestamp 1679581782
transform 1 0 4608 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_49
timestamp 1679581782
transform 1 0 5280 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_56
timestamp 1679581782
transform 1 0 5952 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_63
timestamp 1679581782
transform 1 0 6624 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_70
timestamp 1679581782
transform 1 0 7296 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_77
timestamp 1679581782
transform 1 0 7968 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_84
timestamp 1679581782
transform 1 0 8640 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_91
timestamp 1679581782
transform 1 0 9312 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_98
timestamp 1679581782
transform 1 0 9984 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_105
timestamp 1679581782
transform 1 0 10656 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_112
timestamp 1679581782
transform 1 0 11328 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_119
timestamp 1679581782
transform 1 0 12000 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_126
timestamp 1679581782
transform 1 0 12672 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_133
timestamp 1679581782
transform 1 0 13344 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_140
timestamp 1679581782
transform 1 0 14016 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_4  FILLER_37_147
timestamp 1679577901
transform 1 0 14688 0 -1 29484
box -48 -56 432 834
use sg13g2_fill_2  FILLER_37_151
timestamp 1677580104
transform 1 0 15072 0 -1 29484
box -48 -56 240 834
use sg13g2_decap_8  FILLER_37_180
timestamp 1679581782
transform 1 0 17856 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_187
timestamp 1679581782
transform 1 0 18528 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_194
timestamp 1679581782
transform 1 0 19200 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_201
timestamp 1679581782
transform 1 0 19872 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_208
timestamp 1679581782
transform 1 0 20544 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_215
timestamp 1679581782
transform 1 0 21216 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_222
timestamp 1679581782
transform 1 0 21888 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_229
timestamp 1679581782
transform 1 0 22560 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_236
timestamp 1679581782
transform 1 0 23232 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_243
timestamp 1679581782
transform 1 0 23904 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_250
timestamp 1679581782
transform 1 0 24576 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_257
timestamp 1679581782
transform 1 0 25248 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_264
timestamp 1679581782
transform 1 0 25920 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_271
timestamp 1679581782
transform 1 0 26592 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_278
timestamp 1679581782
transform 1 0 27264 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_285
timestamp 1679581782
transform 1 0 27936 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_292
timestamp 1679581782
transform 1 0 28608 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_299
timestamp 1679581782
transform 1 0 29280 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_306
timestamp 1679581782
transform 1 0 29952 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_4  FILLER_37_313
timestamp 1679577901
transform 1 0 30624 0 -1 29484
box -48 -56 432 834
use sg13g2_fill_1  FILLER_37_317
timestamp 1677579658
transform 1 0 31008 0 -1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_37_321
timestamp 1679581782
transform 1 0 31392 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_328
timestamp 1679581782
transform 1 0 32064 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_335
timestamp 1679581782
transform 1 0 32736 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_342
timestamp 1679581782
transform 1 0 33408 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_349
timestamp 1679581782
transform 1 0 34080 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_356
timestamp 1679581782
transform 1 0 34752 0 -1 29484
box -48 -56 720 834
use sg13g2_fill_1  FILLER_37_363
timestamp 1677579658
transform 1 0 35424 0 -1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_37_370
timestamp 1679581782
transform 1 0 36096 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_377
timestamp 1679581782
transform 1 0 36768 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_384
timestamp 1679581782
transform 1 0 37440 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_391
timestamp 1679581782
transform 1 0 38112 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_398
timestamp 1679581782
transform 1 0 38784 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_405
timestamp 1679581782
transform 1 0 39456 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_412
timestamp 1679581782
transform 1 0 40128 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_419
timestamp 1679581782
transform 1 0 40800 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_426
timestamp 1679581782
transform 1 0 41472 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_433
timestamp 1679581782
transform 1 0 42144 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_440
timestamp 1679581782
transform 1 0 42816 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_447
timestamp 1679581782
transform 1 0 43488 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_454
timestamp 1679581782
transform 1 0 44160 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_461
timestamp 1679581782
transform 1 0 44832 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_468
timestamp 1679581782
transform 1 0 45504 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_475
timestamp 1679581782
transform 1 0 46176 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_482
timestamp 1679581782
transform 1 0 46848 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_489
timestamp 1679581782
transform 1 0 47520 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_496
timestamp 1679581782
transform 1 0 48192 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_503
timestamp 1679581782
transform 1 0 48864 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_510
timestamp 1679581782
transform 1 0 49536 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_517
timestamp 1679581782
transform 1 0 50208 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_524
timestamp 1679581782
transform 1 0 50880 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_531
timestamp 1679581782
transform 1 0 51552 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_538
timestamp 1679581782
transform 1 0 52224 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_545
timestamp 1679581782
transform 1 0 52896 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_552
timestamp 1679581782
transform 1 0 53568 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_559
timestamp 1679581782
transform 1 0 54240 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_566
timestamp 1679581782
transform 1 0 54912 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_573
timestamp 1679581782
transform 1 0 55584 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_580
timestamp 1679581782
transform 1 0 56256 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_587
timestamp 1679581782
transform 1 0 56928 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_594
timestamp 1679581782
transform 1 0 57600 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_601
timestamp 1679581782
transform 1 0 58272 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_608
timestamp 1679581782
transform 1 0 58944 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_615
timestamp 1679581782
transform 1 0 59616 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_622
timestamp 1679581782
transform 1 0 60288 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_629
timestamp 1679581782
transform 1 0 60960 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_636
timestamp 1679581782
transform 1 0 61632 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_643
timestamp 1679581782
transform 1 0 62304 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_650
timestamp 1679581782
transform 1 0 62976 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_657
timestamp 1679581782
transform 1 0 63648 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_664
timestamp 1679581782
transform 1 0 64320 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_671
timestamp 1679581782
transform 1 0 64992 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_678
timestamp 1679581782
transform 1 0 65664 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_685
timestamp 1679581782
transform 1 0 66336 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_692
timestamp 1679581782
transform 1 0 67008 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_699
timestamp 1679581782
transform 1 0 67680 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_706
timestamp 1679581782
transform 1 0 68352 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_713
timestamp 1679581782
transform 1 0 69024 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_720
timestamp 1679581782
transform 1 0 69696 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_727
timestamp 1679581782
transform 1 0 70368 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_734
timestamp 1679581782
transform 1 0 71040 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_741
timestamp 1679581782
transform 1 0 71712 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_748
timestamp 1679581782
transform 1 0 72384 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_755
timestamp 1679581782
transform 1 0 73056 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_762
timestamp 1679581782
transform 1 0 73728 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_769
timestamp 1679581782
transform 1 0 74400 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_776
timestamp 1679581782
transform 1 0 75072 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_783
timestamp 1679581782
transform 1 0 75744 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_790
timestamp 1679581782
transform 1 0 76416 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_797
timestamp 1679581782
transform 1 0 77088 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_804
timestamp 1679581782
transform 1 0 77760 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_811
timestamp 1679581782
transform 1 0 78432 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_818
timestamp 1679581782
transform 1 0 79104 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_825
timestamp 1679581782
transform 1 0 79776 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_832
timestamp 1679581782
transform 1 0 80448 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_839
timestamp 1679581782
transform 1 0 81120 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_846
timestamp 1679581782
transform 1 0 81792 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_853
timestamp 1679581782
transform 1 0 82464 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_860
timestamp 1679581782
transform 1 0 83136 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_867
timestamp 1679581782
transform 1 0 83808 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_874
timestamp 1679581782
transform 1 0 84480 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_881
timestamp 1679581782
transform 1 0 85152 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_888
timestamp 1679581782
transform 1 0 85824 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_895
timestamp 1679581782
transform 1 0 86496 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_902
timestamp 1679581782
transform 1 0 87168 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_909
timestamp 1679581782
transform 1 0 87840 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_916
timestamp 1679581782
transform 1 0 88512 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_923
timestamp 1679581782
transform 1 0 89184 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_930
timestamp 1679581782
transform 1 0 89856 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_937
timestamp 1679581782
transform 1 0 90528 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_944
timestamp 1679581782
transform 1 0 91200 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_951
timestamp 1679581782
transform 1 0 91872 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_958
timestamp 1679581782
transform 1 0 92544 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_965
timestamp 1679581782
transform 1 0 93216 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_972
timestamp 1679581782
transform 1 0 93888 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_979
timestamp 1679581782
transform 1 0 94560 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_986
timestamp 1679581782
transform 1 0 95232 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_993
timestamp 1679581782
transform 1 0 95904 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_1000
timestamp 1679581782
transform 1 0 96576 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_1007
timestamp 1679581782
transform 1 0 97248 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_1014
timestamp 1679581782
transform 1 0 97920 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_1021
timestamp 1679581782
transform 1 0 98592 0 -1 29484
box -48 -56 720 834
use sg13g2_fill_1  FILLER_37_1028
timestamp 1677579658
transform 1 0 99264 0 -1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_38_4
timestamp 1679581782
transform 1 0 960 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_11
timestamp 1679581782
transform 1 0 1632 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_18
timestamp 1679581782
transform 1 0 2304 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_25
timestamp 1679581782
transform 1 0 2976 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_32
timestamp 1679581782
transform 1 0 3648 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_39
timestamp 1679581782
transform 1 0 4320 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_46
timestamp 1679581782
transform 1 0 4992 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_53
timestamp 1679581782
transform 1 0 5664 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_60
timestamp 1679581782
transform 1 0 6336 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_67
timestamp 1679581782
transform 1 0 7008 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_74
timestamp 1679581782
transform 1 0 7680 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_81
timestamp 1679581782
transform 1 0 8352 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_88
timestamp 1679581782
transform 1 0 9024 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_95
timestamp 1679581782
transform 1 0 9696 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_102
timestamp 1679581782
transform 1 0 10368 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_109
timestamp 1679581782
transform 1 0 11040 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_116
timestamp 1679581782
transform 1 0 11712 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_123
timestamp 1679581782
transform 1 0 12384 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_130
timestamp 1679581782
transform 1 0 13056 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_137
timestamp 1679581782
transform 1 0 13728 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_144
timestamp 1679581782
transform 1 0 14400 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_151
timestamp 1679581782
transform 1 0 15072 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_158
timestamp 1679581782
transform 1 0 15744 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_165
timestamp 1679581782
transform 1 0 16416 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_172
timestamp 1679581782
transform 1 0 17088 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_179
timestamp 1679581782
transform 1 0 17760 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_186
timestamp 1679581782
transform 1 0 18432 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_193
timestamp 1679581782
transform 1 0 19104 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_200
timestamp 1679581782
transform 1 0 19776 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_207
timestamp 1679581782
transform 1 0 20448 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_214
timestamp 1679581782
transform 1 0 21120 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_221
timestamp 1679581782
transform 1 0 21792 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_228
timestamp 1679581782
transform 1 0 22464 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_235
timestamp 1679581782
transform 1 0 23136 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_242
timestamp 1679581782
transform 1 0 23808 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_249
timestamp 1679581782
transform 1 0 24480 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_256
timestamp 1679581782
transform 1 0 25152 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_263
timestamp 1679581782
transform 1 0 25824 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_270
timestamp 1679581782
transform 1 0 26496 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_277
timestamp 1679581782
transform 1 0 27168 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_284
timestamp 1679581782
transform 1 0 27840 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_291
timestamp 1679581782
transform 1 0 28512 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_298
timestamp 1679581782
transform 1 0 29184 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_305
timestamp 1679581782
transform 1 0 29856 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_312
timestamp 1679581782
transform 1 0 30528 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_319
timestamp 1679581782
transform 1 0 31200 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_326
timestamp 1679581782
transform 1 0 31872 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_333
timestamp 1679581782
transform 1 0 32544 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_340
timestamp 1679581782
transform 1 0 33216 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_347
timestamp 1679581782
transform 1 0 33888 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_354
timestamp 1679581782
transform 1 0 34560 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_361
timestamp 1679581782
transform 1 0 35232 0 1 29484
box -48 -56 720 834
use sg13g2_decap_4  FILLER_38_368
timestamp 1679577901
transform 1 0 35904 0 1 29484
box -48 -56 432 834
use sg13g2_fill_1  FILLER_38_372
timestamp 1677579658
transform 1 0 36288 0 1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_38_379
timestamp 1679581782
transform 1 0 36960 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_386
timestamp 1679581782
transform 1 0 37632 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_393
timestamp 1679581782
transform 1 0 38304 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_400
timestamp 1679581782
transform 1 0 38976 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_407
timestamp 1679581782
transform 1 0 39648 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_414
timestamp 1679581782
transform 1 0 40320 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_421
timestamp 1679581782
transform 1 0 40992 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_428
timestamp 1679581782
transform 1 0 41664 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_435
timestamp 1679581782
transform 1 0 42336 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_442
timestamp 1679581782
transform 1 0 43008 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_449
timestamp 1679581782
transform 1 0 43680 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_456
timestamp 1679581782
transform 1 0 44352 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_463
timestamp 1679581782
transform 1 0 45024 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_470
timestamp 1679581782
transform 1 0 45696 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_477
timestamp 1679581782
transform 1 0 46368 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_484
timestamp 1679581782
transform 1 0 47040 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_491
timestamp 1679581782
transform 1 0 47712 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_498
timestamp 1679581782
transform 1 0 48384 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_505
timestamp 1679581782
transform 1 0 49056 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_512
timestamp 1679581782
transform 1 0 49728 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_519
timestamp 1679581782
transform 1 0 50400 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_526
timestamp 1679581782
transform 1 0 51072 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_533
timestamp 1679581782
transform 1 0 51744 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_540
timestamp 1679581782
transform 1 0 52416 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_547
timestamp 1679581782
transform 1 0 53088 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_554
timestamp 1679581782
transform 1 0 53760 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_561
timestamp 1679581782
transform 1 0 54432 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_568
timestamp 1679581782
transform 1 0 55104 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_575
timestamp 1679581782
transform 1 0 55776 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_582
timestamp 1679581782
transform 1 0 56448 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_589
timestamp 1679581782
transform 1 0 57120 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_596
timestamp 1679581782
transform 1 0 57792 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_603
timestamp 1679581782
transform 1 0 58464 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_610
timestamp 1679581782
transform 1 0 59136 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_617
timestamp 1679581782
transform 1 0 59808 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_624
timestamp 1679581782
transform 1 0 60480 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_631
timestamp 1679581782
transform 1 0 61152 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_638
timestamp 1679581782
transform 1 0 61824 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_645
timestamp 1679581782
transform 1 0 62496 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_652
timestamp 1679581782
transform 1 0 63168 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_659
timestamp 1679581782
transform 1 0 63840 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_666
timestamp 1679581782
transform 1 0 64512 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_673
timestamp 1679581782
transform 1 0 65184 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_680
timestamp 1679581782
transform 1 0 65856 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_687
timestamp 1679581782
transform 1 0 66528 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_694
timestamp 1679581782
transform 1 0 67200 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_701
timestamp 1679581782
transform 1 0 67872 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_708
timestamp 1679581782
transform 1 0 68544 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_715
timestamp 1679581782
transform 1 0 69216 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_722
timestamp 1679581782
transform 1 0 69888 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_729
timestamp 1679581782
transform 1 0 70560 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_736
timestamp 1679581782
transform 1 0 71232 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_743
timestamp 1679581782
transform 1 0 71904 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_750
timestamp 1679581782
transform 1 0 72576 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_757
timestamp 1679581782
transform 1 0 73248 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_764
timestamp 1679581782
transform 1 0 73920 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_771
timestamp 1679581782
transform 1 0 74592 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_778
timestamp 1679581782
transform 1 0 75264 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_785
timestamp 1679581782
transform 1 0 75936 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_792
timestamp 1679581782
transform 1 0 76608 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_799
timestamp 1679581782
transform 1 0 77280 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_806
timestamp 1679581782
transform 1 0 77952 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_813
timestamp 1679581782
transform 1 0 78624 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_820
timestamp 1679581782
transform 1 0 79296 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_827
timestamp 1679581782
transform 1 0 79968 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_834
timestamp 1679581782
transform 1 0 80640 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_841
timestamp 1679581782
transform 1 0 81312 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_848
timestamp 1679581782
transform 1 0 81984 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_855
timestamp 1679581782
transform 1 0 82656 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_862
timestamp 1679581782
transform 1 0 83328 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_869
timestamp 1679581782
transform 1 0 84000 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_876
timestamp 1679581782
transform 1 0 84672 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_883
timestamp 1679581782
transform 1 0 85344 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_890
timestamp 1679581782
transform 1 0 86016 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_897
timestamp 1679581782
transform 1 0 86688 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_904
timestamp 1679581782
transform 1 0 87360 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_911
timestamp 1679581782
transform 1 0 88032 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_918
timestamp 1679581782
transform 1 0 88704 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_925
timestamp 1679581782
transform 1 0 89376 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_932
timestamp 1679581782
transform 1 0 90048 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_939
timestamp 1679581782
transform 1 0 90720 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_946
timestamp 1679581782
transform 1 0 91392 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_953
timestamp 1679581782
transform 1 0 92064 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_960
timestamp 1679581782
transform 1 0 92736 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_967
timestamp 1679581782
transform 1 0 93408 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_974
timestamp 1679581782
transform 1 0 94080 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_981
timestamp 1679581782
transform 1 0 94752 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_988
timestamp 1679581782
transform 1 0 95424 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_995
timestamp 1679581782
transform 1 0 96096 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_1002
timestamp 1679581782
transform 1 0 96768 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_1009
timestamp 1679581782
transform 1 0 97440 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_1016
timestamp 1679581782
transform 1 0 98112 0 1 29484
box -48 -56 720 834
use sg13g2_decap_4  FILLER_38_1023
timestamp 1679577901
transform 1 0 98784 0 1 29484
box -48 -56 432 834
use sg13g2_fill_2  FILLER_38_1027
timestamp 1677580104
transform 1 0 99168 0 1 29484
box -48 -56 240 834
use sg13g2_decap_8  FILLER_39_4
timestamp 1679581782
transform 1 0 960 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_11
timestamp 1679581782
transform 1 0 1632 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_18
timestamp 1679581782
transform 1 0 2304 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_25
timestamp 1679581782
transform 1 0 2976 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_32
timestamp 1679581782
transform 1 0 3648 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_39
timestamp 1679581782
transform 1 0 4320 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_46
timestamp 1679581782
transform 1 0 4992 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_53
timestamp 1679581782
transform 1 0 5664 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_60
timestamp 1679581782
transform 1 0 6336 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_67
timestamp 1679581782
transform 1 0 7008 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_74
timestamp 1679581782
transform 1 0 7680 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_81
timestamp 1679581782
transform 1 0 8352 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_88
timestamp 1679581782
transform 1 0 9024 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_95
timestamp 1679581782
transform 1 0 9696 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_102
timestamp 1679581782
transform 1 0 10368 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_109
timestamp 1679581782
transform 1 0 11040 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_116
timestamp 1679581782
transform 1 0 11712 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_123
timestamp 1679581782
transform 1 0 12384 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_130
timestamp 1679581782
transform 1 0 13056 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_137
timestamp 1679581782
transform 1 0 13728 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_144
timestamp 1679581782
transform 1 0 14400 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_151
timestamp 1679581782
transform 1 0 15072 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_158
timestamp 1679581782
transform 1 0 15744 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_165
timestamp 1679581782
transform 1 0 16416 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_172
timestamp 1679581782
transform 1 0 17088 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_179
timestamp 1679581782
transform 1 0 17760 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_186
timestamp 1679581782
transform 1 0 18432 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_193
timestamp 1679581782
transform 1 0 19104 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_200
timestamp 1679581782
transform 1 0 19776 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_207
timestamp 1679581782
transform 1 0 20448 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_214
timestamp 1679581782
transform 1 0 21120 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_221
timestamp 1679581782
transform 1 0 21792 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_228
timestamp 1679581782
transform 1 0 22464 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_235
timestamp 1679581782
transform 1 0 23136 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_242
timestamp 1679581782
transform 1 0 23808 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_249
timestamp 1679581782
transform 1 0 24480 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_256
timestamp 1679581782
transform 1 0 25152 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_263
timestamp 1679581782
transform 1 0 25824 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_270
timestamp 1679581782
transform 1 0 26496 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_283
timestamp 1679581782
transform 1 0 27744 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_290
timestamp 1679581782
transform 1 0 28416 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_297
timestamp 1679581782
transform 1 0 29088 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_304
timestamp 1679581782
transform 1 0 29760 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_311
timestamp 1679581782
transform 1 0 30432 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_318
timestamp 1679581782
transform 1 0 31104 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_325
timestamp 1679581782
transform 1 0 31776 0 -1 30996
box -48 -56 720 834
use sg13g2_fill_2  FILLER_39_332
timestamp 1677580104
transform 1 0 32448 0 -1 30996
box -48 -56 240 834
use sg13g2_decap_8  FILLER_39_361
timestamp 1679581782
transform 1 0 35232 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_368
timestamp 1679581782
transform 1 0 35904 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_375
timestamp 1679581782
transform 1 0 36576 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_382
timestamp 1679581782
transform 1 0 37248 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_389
timestamp 1679581782
transform 1 0 37920 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_396
timestamp 1679581782
transform 1 0 38592 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_403
timestamp 1679581782
transform 1 0 39264 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_410
timestamp 1679581782
transform 1 0 39936 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_417
timestamp 1679581782
transform 1 0 40608 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_424
timestamp 1679581782
transform 1 0 41280 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_431
timestamp 1679581782
transform 1 0 41952 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_438
timestamp 1679581782
transform 1 0 42624 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_445
timestamp 1679581782
transform 1 0 43296 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_452
timestamp 1679581782
transform 1 0 43968 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_459
timestamp 1679581782
transform 1 0 44640 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_466
timestamp 1679581782
transform 1 0 45312 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_473
timestamp 1679581782
transform 1 0 45984 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_480
timestamp 1679581782
transform 1 0 46656 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_487
timestamp 1679581782
transform 1 0 47328 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_494
timestamp 1679581782
transform 1 0 48000 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_501
timestamp 1679581782
transform 1 0 48672 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_508
timestamp 1679581782
transform 1 0 49344 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_515
timestamp 1679581782
transform 1 0 50016 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_522
timestamp 1679581782
transform 1 0 50688 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_529
timestamp 1679581782
transform 1 0 51360 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_536
timestamp 1679581782
transform 1 0 52032 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_543
timestamp 1679581782
transform 1 0 52704 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_550
timestamp 1679581782
transform 1 0 53376 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_557
timestamp 1679581782
transform 1 0 54048 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_564
timestamp 1679581782
transform 1 0 54720 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_571
timestamp 1679581782
transform 1 0 55392 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_578
timestamp 1679581782
transform 1 0 56064 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_585
timestamp 1679581782
transform 1 0 56736 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_592
timestamp 1679581782
transform 1 0 57408 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_599
timestamp 1679581782
transform 1 0 58080 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_606
timestamp 1679581782
transform 1 0 58752 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_613
timestamp 1679581782
transform 1 0 59424 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_620
timestamp 1679581782
transform 1 0 60096 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_627
timestamp 1679581782
transform 1 0 60768 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_634
timestamp 1679581782
transform 1 0 61440 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_641
timestamp 1679581782
transform 1 0 62112 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_648
timestamp 1679581782
transform 1 0 62784 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_655
timestamp 1679581782
transform 1 0 63456 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_662
timestamp 1679581782
transform 1 0 64128 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_669
timestamp 1679581782
transform 1 0 64800 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_676
timestamp 1679581782
transform 1 0 65472 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_683
timestamp 1679581782
transform 1 0 66144 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_690
timestamp 1679581782
transform 1 0 66816 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_697
timestamp 1679581782
transform 1 0 67488 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_704
timestamp 1679581782
transform 1 0 68160 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_711
timestamp 1679581782
transform 1 0 68832 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_718
timestamp 1679581782
transform 1 0 69504 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_725
timestamp 1679581782
transform 1 0 70176 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_732
timestamp 1679581782
transform 1 0 70848 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_739
timestamp 1679581782
transform 1 0 71520 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_746
timestamp 1679581782
transform 1 0 72192 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_753
timestamp 1679581782
transform 1 0 72864 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_760
timestamp 1679581782
transform 1 0 73536 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_767
timestamp 1679581782
transform 1 0 74208 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_774
timestamp 1679581782
transform 1 0 74880 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_781
timestamp 1679581782
transform 1 0 75552 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_788
timestamp 1679581782
transform 1 0 76224 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_795
timestamp 1679581782
transform 1 0 76896 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_802
timestamp 1679581782
transform 1 0 77568 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_809
timestamp 1679581782
transform 1 0 78240 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_816
timestamp 1679581782
transform 1 0 78912 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_823
timestamp 1679581782
transform 1 0 79584 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_830
timestamp 1679581782
transform 1 0 80256 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_837
timestamp 1679581782
transform 1 0 80928 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_844
timestamp 1679581782
transform 1 0 81600 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_851
timestamp 1679581782
transform 1 0 82272 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_858
timestamp 1679581782
transform 1 0 82944 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_865
timestamp 1679581782
transform 1 0 83616 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_872
timestamp 1679581782
transform 1 0 84288 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_879
timestamp 1679581782
transform 1 0 84960 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_886
timestamp 1679581782
transform 1 0 85632 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_893
timestamp 1679581782
transform 1 0 86304 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_900
timestamp 1679581782
transform 1 0 86976 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_907
timestamp 1679581782
transform 1 0 87648 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_914
timestamp 1679581782
transform 1 0 88320 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_921
timestamp 1679581782
transform 1 0 88992 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_928
timestamp 1679581782
transform 1 0 89664 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_935
timestamp 1679581782
transform 1 0 90336 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_942
timestamp 1679581782
transform 1 0 91008 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_949
timestamp 1679581782
transform 1 0 91680 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_956
timestamp 1679581782
transform 1 0 92352 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_963
timestamp 1679581782
transform 1 0 93024 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_970
timestamp 1679581782
transform 1 0 93696 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_977
timestamp 1679581782
transform 1 0 94368 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_984
timestamp 1679581782
transform 1 0 95040 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_991
timestamp 1679581782
transform 1 0 95712 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_998
timestamp 1679581782
transform 1 0 96384 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_1005
timestamp 1679581782
transform 1 0 97056 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_1012
timestamp 1679581782
transform 1 0 97728 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_1019
timestamp 1679581782
transform 1 0 98400 0 -1 30996
box -48 -56 720 834
use sg13g2_fill_2  FILLER_39_1026
timestamp 1677580104
transform 1 0 99072 0 -1 30996
box -48 -56 240 834
use sg13g2_fill_1  FILLER_39_1028
timestamp 1677579658
transform 1 0 99264 0 -1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_40_4
timestamp 1679581782
transform 1 0 960 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_11
timestamp 1679581782
transform 1 0 1632 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_18
timestamp 1679581782
transform 1 0 2304 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_25
timestamp 1679581782
transform 1 0 2976 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_32
timestamp 1679581782
transform 1 0 3648 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_39
timestamp 1679581782
transform 1 0 4320 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_46
timestamp 1679581782
transform 1 0 4992 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_53
timestamp 1679581782
transform 1 0 5664 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_60
timestamp 1679581782
transform 1 0 6336 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_67
timestamp 1679581782
transform 1 0 7008 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_74
timestamp 1679581782
transform 1 0 7680 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_81
timestamp 1679581782
transform 1 0 8352 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_88
timestamp 1679581782
transform 1 0 9024 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_95
timestamp 1679581782
transform 1 0 9696 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_102
timestamp 1679581782
transform 1 0 10368 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_109
timestamp 1679581782
transform 1 0 11040 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_116
timestamp 1679581782
transform 1 0 11712 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_123
timestamp 1679581782
transform 1 0 12384 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_130
timestamp 1679581782
transform 1 0 13056 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_137
timestamp 1679581782
transform 1 0 13728 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_144
timestamp 1679581782
transform 1 0 14400 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_151
timestamp 1679581782
transform 1 0 15072 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_158
timestamp 1679581782
transform 1 0 15744 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_165
timestamp 1679581782
transform 1 0 16416 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_172
timestamp 1679581782
transform 1 0 17088 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_179
timestamp 1679581782
transform 1 0 17760 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_186
timestamp 1679581782
transform 1 0 18432 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_193
timestamp 1679581782
transform 1 0 19104 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_200
timestamp 1679581782
transform 1 0 19776 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_207
timestamp 1679581782
transform 1 0 20448 0 1 30996
box -48 -56 720 834
use sg13g2_fill_2  FILLER_40_214
timestamp 1677580104
transform 1 0 21120 0 1 30996
box -48 -56 240 834
use sg13g2_decap_8  FILLER_40_243
timestamp 1679581782
transform 1 0 23904 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_250
timestamp 1679581782
transform 1 0 24576 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_257
timestamp 1679581782
transform 1 0 25248 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_264
timestamp 1679581782
transform 1 0 25920 0 1 30996
box -48 -56 720 834
use sg13g2_fill_1  FILLER_40_271
timestamp 1677579658
transform 1 0 26592 0 1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_40_299
timestamp 1679581782
transform 1 0 29280 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_306
timestamp 1679581782
transform 1 0 29952 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_313
timestamp 1679581782
transform 1 0 30624 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_320
timestamp 1679581782
transform 1 0 31296 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_327
timestamp 1679581782
transform 1 0 31968 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_334
timestamp 1679581782
transform 1 0 32640 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_341
timestamp 1679581782
transform 1 0 33312 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_348
timestamp 1679581782
transform 1 0 33984 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_355
timestamp 1679581782
transform 1 0 34656 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_362
timestamp 1679581782
transform 1 0 35328 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_369
timestamp 1679581782
transform 1 0 36000 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_376
timestamp 1679581782
transform 1 0 36672 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_383
timestamp 1679581782
transform 1 0 37344 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_390
timestamp 1679581782
transform 1 0 38016 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_397
timestamp 1679581782
transform 1 0 38688 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_404
timestamp 1679581782
transform 1 0 39360 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_411
timestamp 1679581782
transform 1 0 40032 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_418
timestamp 1679581782
transform 1 0 40704 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_425
timestamp 1679581782
transform 1 0 41376 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_432
timestamp 1679581782
transform 1 0 42048 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_439
timestamp 1679581782
transform 1 0 42720 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_446
timestamp 1679581782
transform 1 0 43392 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_453
timestamp 1679581782
transform 1 0 44064 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_460
timestamp 1679581782
transform 1 0 44736 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_467
timestamp 1679581782
transform 1 0 45408 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_474
timestamp 1679581782
transform 1 0 46080 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_481
timestamp 1679581782
transform 1 0 46752 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_488
timestamp 1679581782
transform 1 0 47424 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_495
timestamp 1679581782
transform 1 0 48096 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_502
timestamp 1679581782
transform 1 0 48768 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_509
timestamp 1679581782
transform 1 0 49440 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_516
timestamp 1679581782
transform 1 0 50112 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_523
timestamp 1679581782
transform 1 0 50784 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_530
timestamp 1679581782
transform 1 0 51456 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_537
timestamp 1679581782
transform 1 0 52128 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_544
timestamp 1679581782
transform 1 0 52800 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_551
timestamp 1679581782
transform 1 0 53472 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_558
timestamp 1679581782
transform 1 0 54144 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_565
timestamp 1679581782
transform 1 0 54816 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_572
timestamp 1679581782
transform 1 0 55488 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_579
timestamp 1679581782
transform 1 0 56160 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_586
timestamp 1679581782
transform 1 0 56832 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_593
timestamp 1679581782
transform 1 0 57504 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_600
timestamp 1679581782
transform 1 0 58176 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_607
timestamp 1679581782
transform 1 0 58848 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_614
timestamp 1679581782
transform 1 0 59520 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_621
timestamp 1679581782
transform 1 0 60192 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_628
timestamp 1679581782
transform 1 0 60864 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_635
timestamp 1679581782
transform 1 0 61536 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_642
timestamp 1679581782
transform 1 0 62208 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_649
timestamp 1679581782
transform 1 0 62880 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_656
timestamp 1679581782
transform 1 0 63552 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_663
timestamp 1679581782
transform 1 0 64224 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_670
timestamp 1679581782
transform 1 0 64896 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_677
timestamp 1679581782
transform 1 0 65568 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_684
timestamp 1679581782
transform 1 0 66240 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_691
timestamp 1679581782
transform 1 0 66912 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_698
timestamp 1679581782
transform 1 0 67584 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_705
timestamp 1679581782
transform 1 0 68256 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_712
timestamp 1679581782
transform 1 0 68928 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_719
timestamp 1679581782
transform 1 0 69600 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_726
timestamp 1679581782
transform 1 0 70272 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_733
timestamp 1679581782
transform 1 0 70944 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_740
timestamp 1679581782
transform 1 0 71616 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_747
timestamp 1679581782
transform 1 0 72288 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_754
timestamp 1679581782
transform 1 0 72960 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_761
timestamp 1679581782
transform 1 0 73632 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_768
timestamp 1679581782
transform 1 0 74304 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_775
timestamp 1679581782
transform 1 0 74976 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_782
timestamp 1679581782
transform 1 0 75648 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_789
timestamp 1679581782
transform 1 0 76320 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_796
timestamp 1679581782
transform 1 0 76992 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_803
timestamp 1679581782
transform 1 0 77664 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_810
timestamp 1679581782
transform 1 0 78336 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_817
timestamp 1679581782
transform 1 0 79008 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_824
timestamp 1679581782
transform 1 0 79680 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_831
timestamp 1679581782
transform 1 0 80352 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_838
timestamp 1679581782
transform 1 0 81024 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_845
timestamp 1679581782
transform 1 0 81696 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_852
timestamp 1679581782
transform 1 0 82368 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_859
timestamp 1679581782
transform 1 0 83040 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_866
timestamp 1679581782
transform 1 0 83712 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_873
timestamp 1679581782
transform 1 0 84384 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_880
timestamp 1679581782
transform 1 0 85056 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_887
timestamp 1679581782
transform 1 0 85728 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_894
timestamp 1679581782
transform 1 0 86400 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_901
timestamp 1679581782
transform 1 0 87072 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_908
timestamp 1679581782
transform 1 0 87744 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_915
timestamp 1679581782
transform 1 0 88416 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_922
timestamp 1679581782
transform 1 0 89088 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_929
timestamp 1679581782
transform 1 0 89760 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_936
timestamp 1679581782
transform 1 0 90432 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_943
timestamp 1679581782
transform 1 0 91104 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_950
timestamp 1679581782
transform 1 0 91776 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_957
timestamp 1679581782
transform 1 0 92448 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_964
timestamp 1679581782
transform 1 0 93120 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_971
timestamp 1679581782
transform 1 0 93792 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_978
timestamp 1679581782
transform 1 0 94464 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_985
timestamp 1679581782
transform 1 0 95136 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_992
timestamp 1679581782
transform 1 0 95808 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_999
timestamp 1679581782
transform 1 0 96480 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_1006
timestamp 1679581782
transform 1 0 97152 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_1013
timestamp 1679581782
transform 1 0 97824 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_1020
timestamp 1679581782
transform 1 0 98496 0 1 30996
box -48 -56 720 834
use sg13g2_fill_2  FILLER_40_1027
timestamp 1677580104
transform 1 0 99168 0 1 30996
box -48 -56 240 834
use sg13g2_decap_8  FILLER_41_4
timestamp 1679581782
transform 1 0 960 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_11
timestamp 1679581782
transform 1 0 1632 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_18
timestamp 1679581782
transform 1 0 2304 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_25
timestamp 1679581782
transform 1 0 2976 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_32
timestamp 1679581782
transform 1 0 3648 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_39
timestamp 1679581782
transform 1 0 4320 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_46
timestamp 1679581782
transform 1 0 4992 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_53
timestamp 1679581782
transform 1 0 5664 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_60
timestamp 1679581782
transform 1 0 6336 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_67
timestamp 1679581782
transform 1 0 7008 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_74
timestamp 1679581782
transform 1 0 7680 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_81
timestamp 1679581782
transform 1 0 8352 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_88
timestamp 1679581782
transform 1 0 9024 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_95
timestamp 1679581782
transform 1 0 9696 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_102
timestamp 1679581782
transform 1 0 10368 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_109
timestamp 1679581782
transform 1 0 11040 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_116
timestamp 1679581782
transform 1 0 11712 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_123
timestamp 1679581782
transform 1 0 12384 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_130
timestamp 1679581782
transform 1 0 13056 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_137
timestamp 1679581782
transform 1 0 13728 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_144
timestamp 1679581782
transform 1 0 14400 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_151
timestamp 1679581782
transform 1 0 15072 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_158
timestamp 1679581782
transform 1 0 15744 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_165
timestamp 1679581782
transform 1 0 16416 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_172
timestamp 1679581782
transform 1 0 17088 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_179
timestamp 1679581782
transform 1 0 17760 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_186
timestamp 1679581782
transform 1 0 18432 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_193
timestamp 1679581782
transform 1 0 19104 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_200
timestamp 1679581782
transform 1 0 19776 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_207
timestamp 1679581782
transform 1 0 20448 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_214
timestamp 1679581782
transform 1 0 21120 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_221
timestamp 1679581782
transform 1 0 21792 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_228
timestamp 1679581782
transform 1 0 22464 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_235
timestamp 1679581782
transform 1 0 23136 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_242
timestamp 1679581782
transform 1 0 23808 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_249
timestamp 1679581782
transform 1 0 24480 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_256
timestamp 1679581782
transform 1 0 25152 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_263
timestamp 1679581782
transform 1 0 25824 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_270
timestamp 1679581782
transform 1 0 26496 0 -1 32508
box -48 -56 720 834
use sg13g2_fill_2  FILLER_41_277
timestamp 1677580104
transform 1 0 27168 0 -1 32508
box -48 -56 240 834
use sg13g2_decap_8  FILLER_41_285
timestamp 1679581782
transform 1 0 27936 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_292
timestamp 1679581782
transform 1 0 28608 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_299
timestamp 1679581782
transform 1 0 29280 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_306
timestamp 1679581782
transform 1 0 29952 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_313
timestamp 1679581782
transform 1 0 30624 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_320
timestamp 1679581782
transform 1 0 31296 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_327
timestamp 1679581782
transform 1 0 31968 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_334
timestamp 1679581782
transform 1 0 32640 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_341
timestamp 1679581782
transform 1 0 33312 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_348
timestamp 1679581782
transform 1 0 33984 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_355
timestamp 1679581782
transform 1 0 34656 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_362
timestamp 1679581782
transform 1 0 35328 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_369
timestamp 1679581782
transform 1 0 36000 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_376
timestamp 1679581782
transform 1 0 36672 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_383
timestamp 1679581782
transform 1 0 37344 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_390
timestamp 1679581782
transform 1 0 38016 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_397
timestamp 1679581782
transform 1 0 38688 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_404
timestamp 1679581782
transform 1 0 39360 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_411
timestamp 1679581782
transform 1 0 40032 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_418
timestamp 1679581782
transform 1 0 40704 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_425
timestamp 1679581782
transform 1 0 41376 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_432
timestamp 1679581782
transform 1 0 42048 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_439
timestamp 1679581782
transform 1 0 42720 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_446
timestamp 1679581782
transform 1 0 43392 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_453
timestamp 1679581782
transform 1 0 44064 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_460
timestamp 1679581782
transform 1 0 44736 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_467
timestamp 1679581782
transform 1 0 45408 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_474
timestamp 1679581782
transform 1 0 46080 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_481
timestamp 1679581782
transform 1 0 46752 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_488
timestamp 1679581782
transform 1 0 47424 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_495
timestamp 1679581782
transform 1 0 48096 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_502
timestamp 1679581782
transform 1 0 48768 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_509
timestamp 1679581782
transform 1 0 49440 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_516
timestamp 1679581782
transform 1 0 50112 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_523
timestamp 1679581782
transform 1 0 50784 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_530
timestamp 1679581782
transform 1 0 51456 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_537
timestamp 1679581782
transform 1 0 52128 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_544
timestamp 1679581782
transform 1 0 52800 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_551
timestamp 1679581782
transform 1 0 53472 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_558
timestamp 1679581782
transform 1 0 54144 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_565
timestamp 1679581782
transform 1 0 54816 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_572
timestamp 1679581782
transform 1 0 55488 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_579
timestamp 1679581782
transform 1 0 56160 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_586
timestamp 1679581782
transform 1 0 56832 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_593
timestamp 1679581782
transform 1 0 57504 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_600
timestamp 1679581782
transform 1 0 58176 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_607
timestamp 1679581782
transform 1 0 58848 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_614
timestamp 1679581782
transform 1 0 59520 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_621
timestamp 1679581782
transform 1 0 60192 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_628
timestamp 1679581782
transform 1 0 60864 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_635
timestamp 1679581782
transform 1 0 61536 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_642
timestamp 1679581782
transform 1 0 62208 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_649
timestamp 1679581782
transform 1 0 62880 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_656
timestamp 1679581782
transform 1 0 63552 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_663
timestamp 1679581782
transform 1 0 64224 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_670
timestamp 1679581782
transform 1 0 64896 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_677
timestamp 1679581782
transform 1 0 65568 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_684
timestamp 1679581782
transform 1 0 66240 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_691
timestamp 1679581782
transform 1 0 66912 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_698
timestamp 1679581782
transform 1 0 67584 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_705
timestamp 1679581782
transform 1 0 68256 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_712
timestamp 1679581782
transform 1 0 68928 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_719
timestamp 1679581782
transform 1 0 69600 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_726
timestamp 1679581782
transform 1 0 70272 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_733
timestamp 1679581782
transform 1 0 70944 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_740
timestamp 1679581782
transform 1 0 71616 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_747
timestamp 1679581782
transform 1 0 72288 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_754
timestamp 1679581782
transform 1 0 72960 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_761
timestamp 1679581782
transform 1 0 73632 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_768
timestamp 1679581782
transform 1 0 74304 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_775
timestamp 1679581782
transform 1 0 74976 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_782
timestamp 1679581782
transform 1 0 75648 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_789
timestamp 1679581782
transform 1 0 76320 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_796
timestamp 1679581782
transform 1 0 76992 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_803
timestamp 1679581782
transform 1 0 77664 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_810
timestamp 1679581782
transform 1 0 78336 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_817
timestamp 1679581782
transform 1 0 79008 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_824
timestamp 1679581782
transform 1 0 79680 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_831
timestamp 1679581782
transform 1 0 80352 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_838
timestamp 1679581782
transform 1 0 81024 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_845
timestamp 1679581782
transform 1 0 81696 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_852
timestamp 1679581782
transform 1 0 82368 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_859
timestamp 1679581782
transform 1 0 83040 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_866
timestamp 1679581782
transform 1 0 83712 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_873
timestamp 1679581782
transform 1 0 84384 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_880
timestamp 1679581782
transform 1 0 85056 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_887
timestamp 1679581782
transform 1 0 85728 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_894
timestamp 1679581782
transform 1 0 86400 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_901
timestamp 1679581782
transform 1 0 87072 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_908
timestamp 1679581782
transform 1 0 87744 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_915
timestamp 1679581782
transform 1 0 88416 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_922
timestamp 1679581782
transform 1 0 89088 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_929
timestamp 1679581782
transform 1 0 89760 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_936
timestamp 1679581782
transform 1 0 90432 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_943
timestamp 1679581782
transform 1 0 91104 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_950
timestamp 1679581782
transform 1 0 91776 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_957
timestamp 1679581782
transform 1 0 92448 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_964
timestamp 1679581782
transform 1 0 93120 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_971
timestamp 1679581782
transform 1 0 93792 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_978
timestamp 1679581782
transform 1 0 94464 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_985
timestamp 1679581782
transform 1 0 95136 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_992
timestamp 1679581782
transform 1 0 95808 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_999
timestamp 1679581782
transform 1 0 96480 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_1006
timestamp 1679581782
transform 1 0 97152 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_1013
timestamp 1679581782
transform 1 0 97824 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_1020
timestamp 1679581782
transform 1 0 98496 0 -1 32508
box -48 -56 720 834
use sg13g2_fill_2  FILLER_41_1027
timestamp 1677580104
transform 1 0 99168 0 -1 32508
box -48 -56 240 834
use sg13g2_decap_8  FILLER_42_5
timestamp 1679581782
transform 1 0 1056 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_12
timestamp 1679581782
transform 1 0 1728 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_19
timestamp 1679581782
transform 1 0 2400 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_26
timestamp 1679581782
transform 1 0 3072 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_33
timestamp 1679581782
transform 1 0 3744 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_40
timestamp 1679581782
transform 1 0 4416 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_47
timestamp 1679581782
transform 1 0 5088 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_54
timestamp 1679581782
transform 1 0 5760 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_61
timestamp 1679581782
transform 1 0 6432 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_68
timestamp 1679581782
transform 1 0 7104 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_75
timestamp 1679581782
transform 1 0 7776 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_82
timestamp 1679581782
transform 1 0 8448 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_89
timestamp 1679581782
transform 1 0 9120 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_96
timestamp 1679581782
transform 1 0 9792 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_103
timestamp 1679581782
transform 1 0 10464 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_110
timestamp 1679581782
transform 1 0 11136 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_117
timestamp 1679581782
transform 1 0 11808 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_124
timestamp 1679581782
transform 1 0 12480 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_131
timestamp 1679581782
transform 1 0 13152 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_138
timestamp 1679581782
transform 1 0 13824 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_145
timestamp 1679581782
transform 1 0 14496 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_152
timestamp 1679581782
transform 1 0 15168 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_159
timestamp 1679581782
transform 1 0 15840 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_166
timestamp 1679581782
transform 1 0 16512 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_173
timestamp 1679581782
transform 1 0 17184 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_180
timestamp 1679581782
transform 1 0 17856 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_187
timestamp 1679581782
transform 1 0 18528 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_194
timestamp 1679581782
transform 1 0 19200 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_201
timestamp 1679581782
transform 1 0 19872 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_208
timestamp 1679581782
transform 1 0 20544 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_215
timestamp 1679581782
transform 1 0 21216 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_222
timestamp 1679581782
transform 1 0 21888 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_229
timestamp 1679581782
transform 1 0 22560 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_236
timestamp 1679581782
transform 1 0 23232 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_243
timestamp 1679581782
transform 1 0 23904 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_250
timestamp 1679581782
transform 1 0 24576 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_257
timestamp 1679581782
transform 1 0 25248 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_264
timestamp 1679581782
transform 1 0 25920 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_271
timestamp 1679581782
transform 1 0 26592 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_278
timestamp 1679581782
transform 1 0 27264 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_285
timestamp 1679581782
transform 1 0 27936 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_292
timestamp 1679581782
transform 1 0 28608 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_299
timestamp 1679581782
transform 1 0 29280 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_306
timestamp 1679581782
transform 1 0 29952 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_313
timestamp 1679581782
transform 1 0 30624 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_320
timestamp 1679581782
transform 1 0 31296 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_327
timestamp 1679581782
transform 1 0 31968 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_334
timestamp 1679581782
transform 1 0 32640 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_341
timestamp 1679581782
transform 1 0 33312 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_348
timestamp 1679581782
transform 1 0 33984 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_355
timestamp 1679581782
transform 1 0 34656 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_362
timestamp 1679581782
transform 1 0 35328 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_369
timestamp 1679581782
transform 1 0 36000 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_376
timestamp 1679581782
transform 1 0 36672 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_383
timestamp 1679581782
transform 1 0 37344 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_390
timestamp 1679581782
transform 1 0 38016 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_397
timestamp 1679581782
transform 1 0 38688 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_404
timestamp 1679581782
transform 1 0 39360 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_411
timestamp 1679581782
transform 1 0 40032 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_418
timestamp 1679581782
transform 1 0 40704 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_425
timestamp 1679581782
transform 1 0 41376 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_432
timestamp 1679581782
transform 1 0 42048 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_439
timestamp 1679581782
transform 1 0 42720 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_446
timestamp 1679581782
transform 1 0 43392 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_453
timestamp 1679581782
transform 1 0 44064 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_460
timestamp 1679581782
transform 1 0 44736 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_467
timestamp 1679581782
transform 1 0 45408 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_474
timestamp 1679581782
transform 1 0 46080 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_481
timestamp 1679581782
transform 1 0 46752 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_488
timestamp 1679581782
transform 1 0 47424 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_495
timestamp 1679581782
transform 1 0 48096 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_502
timestamp 1679581782
transform 1 0 48768 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_509
timestamp 1679581782
transform 1 0 49440 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_516
timestamp 1679581782
transform 1 0 50112 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_523
timestamp 1679581782
transform 1 0 50784 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_530
timestamp 1679581782
transform 1 0 51456 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_537
timestamp 1679581782
transform 1 0 52128 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_544
timestamp 1679581782
transform 1 0 52800 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_551
timestamp 1679581782
transform 1 0 53472 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_558
timestamp 1679581782
transform 1 0 54144 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_565
timestamp 1679581782
transform 1 0 54816 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_572
timestamp 1679581782
transform 1 0 55488 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_579
timestamp 1679581782
transform 1 0 56160 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_586
timestamp 1679581782
transform 1 0 56832 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_593
timestamp 1679581782
transform 1 0 57504 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_600
timestamp 1679581782
transform 1 0 58176 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_607
timestamp 1679581782
transform 1 0 58848 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_614
timestamp 1679581782
transform 1 0 59520 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_621
timestamp 1679581782
transform 1 0 60192 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_628
timestamp 1679581782
transform 1 0 60864 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_635
timestamp 1679581782
transform 1 0 61536 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_642
timestamp 1679581782
transform 1 0 62208 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_649
timestamp 1679581782
transform 1 0 62880 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_656
timestamp 1679581782
transform 1 0 63552 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_663
timestamp 1679581782
transform 1 0 64224 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_670
timestamp 1679581782
transform 1 0 64896 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_677
timestamp 1679581782
transform 1 0 65568 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_684
timestamp 1679581782
transform 1 0 66240 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_691
timestamp 1679581782
transform 1 0 66912 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_698
timestamp 1679581782
transform 1 0 67584 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_705
timestamp 1679581782
transform 1 0 68256 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_712
timestamp 1679581782
transform 1 0 68928 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_719
timestamp 1679581782
transform 1 0 69600 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_726
timestamp 1679581782
transform 1 0 70272 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_733
timestamp 1679581782
transform 1 0 70944 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_740
timestamp 1679581782
transform 1 0 71616 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_747
timestamp 1679581782
transform 1 0 72288 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_754
timestamp 1679581782
transform 1 0 72960 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_761
timestamp 1679581782
transform 1 0 73632 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_768
timestamp 1679581782
transform 1 0 74304 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_775
timestamp 1679581782
transform 1 0 74976 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_782
timestamp 1679581782
transform 1 0 75648 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_789
timestamp 1679581782
transform 1 0 76320 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_796
timestamp 1679581782
transform 1 0 76992 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_803
timestamp 1679581782
transform 1 0 77664 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_810
timestamp 1679581782
transform 1 0 78336 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_817
timestamp 1679581782
transform 1 0 79008 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_824
timestamp 1679581782
transform 1 0 79680 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_831
timestamp 1679581782
transform 1 0 80352 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_838
timestamp 1679581782
transform 1 0 81024 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_845
timestamp 1679581782
transform 1 0 81696 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_852
timestamp 1679581782
transform 1 0 82368 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_859
timestamp 1679581782
transform 1 0 83040 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_866
timestamp 1679581782
transform 1 0 83712 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_873
timestamp 1679581782
transform 1 0 84384 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_880
timestamp 1679581782
transform 1 0 85056 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_887
timestamp 1679581782
transform 1 0 85728 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_894
timestamp 1679581782
transform 1 0 86400 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_901
timestamp 1679581782
transform 1 0 87072 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_908
timestamp 1679581782
transform 1 0 87744 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_915
timestamp 1679581782
transform 1 0 88416 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_922
timestamp 1679581782
transform 1 0 89088 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_929
timestamp 1679581782
transform 1 0 89760 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_936
timestamp 1679581782
transform 1 0 90432 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_943
timestamp 1679581782
transform 1 0 91104 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_950
timestamp 1679581782
transform 1 0 91776 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_957
timestamp 1679581782
transform 1 0 92448 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_964
timestamp 1679581782
transform 1 0 93120 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_971
timestamp 1679581782
transform 1 0 93792 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_978
timestamp 1679581782
transform 1 0 94464 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_985
timestamp 1679581782
transform 1 0 95136 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_992
timestamp 1679581782
transform 1 0 95808 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_999
timestamp 1679581782
transform 1 0 96480 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_1006
timestamp 1679581782
transform 1 0 97152 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_1013
timestamp 1679581782
transform 1 0 97824 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_1020
timestamp 1679581782
transform 1 0 98496 0 1 32508
box -48 -56 720 834
use sg13g2_fill_2  FILLER_42_1027
timestamp 1677580104
transform 1 0 99168 0 1 32508
box -48 -56 240 834
use sg13g2_decap_8  FILLER_43_5
timestamp 1679581782
transform 1 0 1056 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_12
timestamp 1679581782
transform 1 0 1728 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_19
timestamp 1679581782
transform 1 0 2400 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_26
timestamp 1679581782
transform 1 0 3072 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_33
timestamp 1679581782
transform 1 0 3744 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_40
timestamp 1679581782
transform 1 0 4416 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_47
timestamp 1679581782
transform 1 0 5088 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_54
timestamp 1679581782
transform 1 0 5760 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_61
timestamp 1679581782
transform 1 0 6432 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_68
timestamp 1679581782
transform 1 0 7104 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_75
timestamp 1679581782
transform 1 0 7776 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_82
timestamp 1679581782
transform 1 0 8448 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_89
timestamp 1679581782
transform 1 0 9120 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_96
timestamp 1679581782
transform 1 0 9792 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_103
timestamp 1679581782
transform 1 0 10464 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_110
timestamp 1679581782
transform 1 0 11136 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_117
timestamp 1679581782
transform 1 0 11808 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_124
timestamp 1679581782
transform 1 0 12480 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_131
timestamp 1679581782
transform 1 0 13152 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_138
timestamp 1679581782
transform 1 0 13824 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_145
timestamp 1679581782
transform 1 0 14496 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_152
timestamp 1679581782
transform 1 0 15168 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_159
timestamp 1679581782
transform 1 0 15840 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_166
timestamp 1679581782
transform 1 0 16512 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_173
timestamp 1679581782
transform 1 0 17184 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_180
timestamp 1679581782
transform 1 0 17856 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_187
timestamp 1679581782
transform 1 0 18528 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_194
timestamp 1679581782
transform 1 0 19200 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_201
timestamp 1679581782
transform 1 0 19872 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_208
timestamp 1679581782
transform 1 0 20544 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_215
timestamp 1679581782
transform 1 0 21216 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_222
timestamp 1679581782
transform 1 0 21888 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_229
timestamp 1679581782
transform 1 0 22560 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_236
timestamp 1679581782
transform 1 0 23232 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_243
timestamp 1679581782
transform 1 0 23904 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_250
timestamp 1679581782
transform 1 0 24576 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_257
timestamp 1679581782
transform 1 0 25248 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_264
timestamp 1679581782
transform 1 0 25920 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_271
timestamp 1679581782
transform 1 0 26592 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_278
timestamp 1679581782
transform 1 0 27264 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_285
timestamp 1679581782
transform 1 0 27936 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_292
timestamp 1679581782
transform 1 0 28608 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_299
timestamp 1679581782
transform 1 0 29280 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_306
timestamp 1679581782
transform 1 0 29952 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_313
timestamp 1679581782
transform 1 0 30624 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_320
timestamp 1679581782
transform 1 0 31296 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_327
timestamp 1679581782
transform 1 0 31968 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_334
timestamp 1679581782
transform 1 0 32640 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_341
timestamp 1679581782
transform 1 0 33312 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_348
timestamp 1679581782
transform 1 0 33984 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_355
timestamp 1679581782
transform 1 0 34656 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_362
timestamp 1679581782
transform 1 0 35328 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_369
timestamp 1679581782
transform 1 0 36000 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_376
timestamp 1679581782
transform 1 0 36672 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_383
timestamp 1679581782
transform 1 0 37344 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_390
timestamp 1679581782
transform 1 0 38016 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_397
timestamp 1679581782
transform 1 0 38688 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_404
timestamp 1679581782
transform 1 0 39360 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_411
timestamp 1679581782
transform 1 0 40032 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_418
timestamp 1679581782
transform 1 0 40704 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_425
timestamp 1679581782
transform 1 0 41376 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_432
timestamp 1679581782
transform 1 0 42048 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_439
timestamp 1679581782
transform 1 0 42720 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_446
timestamp 1679581782
transform 1 0 43392 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_453
timestamp 1679581782
transform 1 0 44064 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_460
timestamp 1679581782
transform 1 0 44736 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_467
timestamp 1679581782
transform 1 0 45408 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_474
timestamp 1679581782
transform 1 0 46080 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_481
timestamp 1679581782
transform 1 0 46752 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_488
timestamp 1679581782
transform 1 0 47424 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_495
timestamp 1679581782
transform 1 0 48096 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_502
timestamp 1679581782
transform 1 0 48768 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_509
timestamp 1679581782
transform 1 0 49440 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_516
timestamp 1679581782
transform 1 0 50112 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_523
timestamp 1679581782
transform 1 0 50784 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_530
timestamp 1679581782
transform 1 0 51456 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_537
timestamp 1679581782
transform 1 0 52128 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_544
timestamp 1679581782
transform 1 0 52800 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_551
timestamp 1679581782
transform 1 0 53472 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_558
timestamp 1679581782
transform 1 0 54144 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_565
timestamp 1679581782
transform 1 0 54816 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_572
timestamp 1679581782
transform 1 0 55488 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_579
timestamp 1679581782
transform 1 0 56160 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_586
timestamp 1679581782
transform 1 0 56832 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_593
timestamp 1679581782
transform 1 0 57504 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_600
timestamp 1679581782
transform 1 0 58176 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_607
timestamp 1679581782
transform 1 0 58848 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_614
timestamp 1679581782
transform 1 0 59520 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_621
timestamp 1679581782
transform 1 0 60192 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_628
timestamp 1679581782
transform 1 0 60864 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_635
timestamp 1679581782
transform 1 0 61536 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_642
timestamp 1679581782
transform 1 0 62208 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_649
timestamp 1679581782
transform 1 0 62880 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_656
timestamp 1679581782
transform 1 0 63552 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_663
timestamp 1679581782
transform 1 0 64224 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_670
timestamp 1679581782
transform 1 0 64896 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_677
timestamp 1679581782
transform 1 0 65568 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_684
timestamp 1679581782
transform 1 0 66240 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_691
timestamp 1679581782
transform 1 0 66912 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_698
timestamp 1679581782
transform 1 0 67584 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_705
timestamp 1679581782
transform 1 0 68256 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_712
timestamp 1679581782
transform 1 0 68928 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_719
timestamp 1679581782
transform 1 0 69600 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_726
timestamp 1679581782
transform 1 0 70272 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_733
timestamp 1679581782
transform 1 0 70944 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_740
timestamp 1679581782
transform 1 0 71616 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_747
timestamp 1679581782
transform 1 0 72288 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_754
timestamp 1679581782
transform 1 0 72960 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_761
timestamp 1679581782
transform 1 0 73632 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_768
timestamp 1679581782
transform 1 0 74304 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_775
timestamp 1679581782
transform 1 0 74976 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_782
timestamp 1679581782
transform 1 0 75648 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_789
timestamp 1679581782
transform 1 0 76320 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_796
timestamp 1679581782
transform 1 0 76992 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_803
timestamp 1679581782
transform 1 0 77664 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_810
timestamp 1679581782
transform 1 0 78336 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_817
timestamp 1679581782
transform 1 0 79008 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_824
timestamp 1679581782
transform 1 0 79680 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_831
timestamp 1679581782
transform 1 0 80352 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_838
timestamp 1679581782
transform 1 0 81024 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_845
timestamp 1679581782
transform 1 0 81696 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_852
timestamp 1679581782
transform 1 0 82368 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_859
timestamp 1679581782
transform 1 0 83040 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_866
timestamp 1679581782
transform 1 0 83712 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_873
timestamp 1679581782
transform 1 0 84384 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_880
timestamp 1679581782
transform 1 0 85056 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_887
timestamp 1679581782
transform 1 0 85728 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_894
timestamp 1679581782
transform 1 0 86400 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_901
timestamp 1679581782
transform 1 0 87072 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_908
timestamp 1679581782
transform 1 0 87744 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_915
timestamp 1679581782
transform 1 0 88416 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_922
timestamp 1679581782
transform 1 0 89088 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_929
timestamp 1679581782
transform 1 0 89760 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_936
timestamp 1679581782
transform 1 0 90432 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_943
timestamp 1679581782
transform 1 0 91104 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_950
timestamp 1679581782
transform 1 0 91776 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_957
timestamp 1679581782
transform 1 0 92448 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_964
timestamp 1679581782
transform 1 0 93120 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_971
timestamp 1679581782
transform 1 0 93792 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_978
timestamp 1679581782
transform 1 0 94464 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_985
timestamp 1679581782
transform 1 0 95136 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_992
timestamp 1679581782
transform 1 0 95808 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_999
timestamp 1679581782
transform 1 0 96480 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_1006
timestamp 1679581782
transform 1 0 97152 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_1013
timestamp 1679581782
transform 1 0 97824 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_1020
timestamp 1679581782
transform 1 0 98496 0 -1 34020
box -48 -56 720 834
use sg13g2_fill_2  FILLER_43_1027
timestamp 1677580104
transform 1 0 99168 0 -1 34020
box -48 -56 240 834
use sg13g2_decap_8  FILLER_44_5
timestamp 1679581782
transform 1 0 1056 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_12
timestamp 1679581782
transform 1 0 1728 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_19
timestamp 1679581782
transform 1 0 2400 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_26
timestamp 1679581782
transform 1 0 3072 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_33
timestamp 1679581782
transform 1 0 3744 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_40
timestamp 1679581782
transform 1 0 4416 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_47
timestamp 1679581782
transform 1 0 5088 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_54
timestamp 1679581782
transform 1 0 5760 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_61
timestamp 1679581782
transform 1 0 6432 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_68
timestamp 1679581782
transform 1 0 7104 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_75
timestamp 1679581782
transform 1 0 7776 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_82
timestamp 1679581782
transform 1 0 8448 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_89
timestamp 1679581782
transform 1 0 9120 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_96
timestamp 1679581782
transform 1 0 9792 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_103
timestamp 1679581782
transform 1 0 10464 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_110
timestamp 1679581782
transform 1 0 11136 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_117
timestamp 1679581782
transform 1 0 11808 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_124
timestamp 1679581782
transform 1 0 12480 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_131
timestamp 1679581782
transform 1 0 13152 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_138
timestamp 1679581782
transform 1 0 13824 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_145
timestamp 1679581782
transform 1 0 14496 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_152
timestamp 1679581782
transform 1 0 15168 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_159
timestamp 1679581782
transform 1 0 15840 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_166
timestamp 1679581782
transform 1 0 16512 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_173
timestamp 1679581782
transform 1 0 17184 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_180
timestamp 1679581782
transform 1 0 17856 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_187
timestamp 1679581782
transform 1 0 18528 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_194
timestamp 1679581782
transform 1 0 19200 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_201
timestamp 1679581782
transform 1 0 19872 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_208
timestamp 1679581782
transform 1 0 20544 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_215
timestamp 1679581782
transform 1 0 21216 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_222
timestamp 1679581782
transform 1 0 21888 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_229
timestamp 1679581782
transform 1 0 22560 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_236
timestamp 1679581782
transform 1 0 23232 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_243
timestamp 1679581782
transform 1 0 23904 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_250
timestamp 1679581782
transform 1 0 24576 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_257
timestamp 1679581782
transform 1 0 25248 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_264
timestamp 1679581782
transform 1 0 25920 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_271
timestamp 1679581782
transform 1 0 26592 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_278
timestamp 1679581782
transform 1 0 27264 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_285
timestamp 1679581782
transform 1 0 27936 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_292
timestamp 1679581782
transform 1 0 28608 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_299
timestamp 1679581782
transform 1 0 29280 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_306
timestamp 1679581782
transform 1 0 29952 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_313
timestamp 1679581782
transform 1 0 30624 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_320
timestamp 1679581782
transform 1 0 31296 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_327
timestamp 1679581782
transform 1 0 31968 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_334
timestamp 1679581782
transform 1 0 32640 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_341
timestamp 1679581782
transform 1 0 33312 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_348
timestamp 1679581782
transform 1 0 33984 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_355
timestamp 1679581782
transform 1 0 34656 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_362
timestamp 1679581782
transform 1 0 35328 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_369
timestamp 1679581782
transform 1 0 36000 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_376
timestamp 1679581782
transform 1 0 36672 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_383
timestamp 1679581782
transform 1 0 37344 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_390
timestamp 1679581782
transform 1 0 38016 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_397
timestamp 1679581782
transform 1 0 38688 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_404
timestamp 1679581782
transform 1 0 39360 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_411
timestamp 1679581782
transform 1 0 40032 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_418
timestamp 1679581782
transform 1 0 40704 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_425
timestamp 1679581782
transform 1 0 41376 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_432
timestamp 1679581782
transform 1 0 42048 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_439
timestamp 1679581782
transform 1 0 42720 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_446
timestamp 1679581782
transform 1 0 43392 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_453
timestamp 1679581782
transform 1 0 44064 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_460
timestamp 1679581782
transform 1 0 44736 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_467
timestamp 1679581782
transform 1 0 45408 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_474
timestamp 1679581782
transform 1 0 46080 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_481
timestamp 1679581782
transform 1 0 46752 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_488
timestamp 1679581782
transform 1 0 47424 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_495
timestamp 1679581782
transform 1 0 48096 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_502
timestamp 1679581782
transform 1 0 48768 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_509
timestamp 1679581782
transform 1 0 49440 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_516
timestamp 1679581782
transform 1 0 50112 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_523
timestamp 1679581782
transform 1 0 50784 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_530
timestamp 1679581782
transform 1 0 51456 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_537
timestamp 1679581782
transform 1 0 52128 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_544
timestamp 1679581782
transform 1 0 52800 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_551
timestamp 1679581782
transform 1 0 53472 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_558
timestamp 1679581782
transform 1 0 54144 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_565
timestamp 1679581782
transform 1 0 54816 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_572
timestamp 1679581782
transform 1 0 55488 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_579
timestamp 1679581782
transform 1 0 56160 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_586
timestamp 1679581782
transform 1 0 56832 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_593
timestamp 1679581782
transform 1 0 57504 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_600
timestamp 1679581782
transform 1 0 58176 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_607
timestamp 1679581782
transform 1 0 58848 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_614
timestamp 1679581782
transform 1 0 59520 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_621
timestamp 1679581782
transform 1 0 60192 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_628
timestamp 1679581782
transform 1 0 60864 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_635
timestamp 1679581782
transform 1 0 61536 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_642
timestamp 1679581782
transform 1 0 62208 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_649
timestamp 1679581782
transform 1 0 62880 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_656
timestamp 1679581782
transform 1 0 63552 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_663
timestamp 1679581782
transform 1 0 64224 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_670
timestamp 1679581782
transform 1 0 64896 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_677
timestamp 1679581782
transform 1 0 65568 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_684
timestamp 1679581782
transform 1 0 66240 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_691
timestamp 1679581782
transform 1 0 66912 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_698
timestamp 1679581782
transform 1 0 67584 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_705
timestamp 1679581782
transform 1 0 68256 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_712
timestamp 1679581782
transform 1 0 68928 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_719
timestamp 1679581782
transform 1 0 69600 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_726
timestamp 1679581782
transform 1 0 70272 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_733
timestamp 1679581782
transform 1 0 70944 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_740
timestamp 1679581782
transform 1 0 71616 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_747
timestamp 1679581782
transform 1 0 72288 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_754
timestamp 1679581782
transform 1 0 72960 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_761
timestamp 1679581782
transform 1 0 73632 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_768
timestamp 1679581782
transform 1 0 74304 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_775
timestamp 1679581782
transform 1 0 74976 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_782
timestamp 1679581782
transform 1 0 75648 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_789
timestamp 1679581782
transform 1 0 76320 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_796
timestamp 1679581782
transform 1 0 76992 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_803
timestamp 1679581782
transform 1 0 77664 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_810
timestamp 1679581782
transform 1 0 78336 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_817
timestamp 1679581782
transform 1 0 79008 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_824
timestamp 1679581782
transform 1 0 79680 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_831
timestamp 1679581782
transform 1 0 80352 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_838
timestamp 1679581782
transform 1 0 81024 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_845
timestamp 1679581782
transform 1 0 81696 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_852
timestamp 1679581782
transform 1 0 82368 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_859
timestamp 1679581782
transform 1 0 83040 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_866
timestamp 1679581782
transform 1 0 83712 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_873
timestamp 1679581782
transform 1 0 84384 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_880
timestamp 1679581782
transform 1 0 85056 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_887
timestamp 1679581782
transform 1 0 85728 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_894
timestamp 1679581782
transform 1 0 86400 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_901
timestamp 1679581782
transform 1 0 87072 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_908
timestamp 1679581782
transform 1 0 87744 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_915
timestamp 1679581782
transform 1 0 88416 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_922
timestamp 1679581782
transform 1 0 89088 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_929
timestamp 1679581782
transform 1 0 89760 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_936
timestamp 1679581782
transform 1 0 90432 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_943
timestamp 1679581782
transform 1 0 91104 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_950
timestamp 1679581782
transform 1 0 91776 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_957
timestamp 1679581782
transform 1 0 92448 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_964
timestamp 1679581782
transform 1 0 93120 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_971
timestamp 1679581782
transform 1 0 93792 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_978
timestamp 1679581782
transform 1 0 94464 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_985
timestamp 1679581782
transform 1 0 95136 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_992
timestamp 1679581782
transform 1 0 95808 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_999
timestamp 1679581782
transform 1 0 96480 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_1006
timestamp 1679581782
transform 1 0 97152 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_1013
timestamp 1679581782
transform 1 0 97824 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_1020
timestamp 1679581782
transform 1 0 98496 0 1 34020
box -48 -56 720 834
use sg13g2_fill_2  FILLER_44_1027
timestamp 1677580104
transform 1 0 99168 0 1 34020
box -48 -56 240 834
use sg13g2_decap_8  FILLER_45_5
timestamp 1679581782
transform 1 0 1056 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_12
timestamp 1679581782
transform 1 0 1728 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_19
timestamp 1679581782
transform 1 0 2400 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_26
timestamp 1679581782
transform 1 0 3072 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_33
timestamp 1679581782
transform 1 0 3744 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_40
timestamp 1679581782
transform 1 0 4416 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_47
timestamp 1679581782
transform 1 0 5088 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_54
timestamp 1679581782
transform 1 0 5760 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_61
timestamp 1679581782
transform 1 0 6432 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_68
timestamp 1679581782
transform 1 0 7104 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_75
timestamp 1679581782
transform 1 0 7776 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_82
timestamp 1679581782
transform 1 0 8448 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_89
timestamp 1679581782
transform 1 0 9120 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_96
timestamp 1679581782
transform 1 0 9792 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_103
timestamp 1679581782
transform 1 0 10464 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_110
timestamp 1679581782
transform 1 0 11136 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_117
timestamp 1679581782
transform 1 0 11808 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_124
timestamp 1679581782
transform 1 0 12480 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_131
timestamp 1679581782
transform 1 0 13152 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_138
timestamp 1679581782
transform 1 0 13824 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_145
timestamp 1679581782
transform 1 0 14496 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_152
timestamp 1679581782
transform 1 0 15168 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_159
timestamp 1679581782
transform 1 0 15840 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_166
timestamp 1679581782
transform 1 0 16512 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_173
timestamp 1679581782
transform 1 0 17184 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_180
timestamp 1679581782
transform 1 0 17856 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_187
timestamp 1679581782
transform 1 0 18528 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_194
timestamp 1679581782
transform 1 0 19200 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_201
timestamp 1679581782
transform 1 0 19872 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_208
timestamp 1679581782
transform 1 0 20544 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_215
timestamp 1679581782
transform 1 0 21216 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_222
timestamp 1679581782
transform 1 0 21888 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_229
timestamp 1679581782
transform 1 0 22560 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_236
timestamp 1679581782
transform 1 0 23232 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_243
timestamp 1679581782
transform 1 0 23904 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_250
timestamp 1679581782
transform 1 0 24576 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_257
timestamp 1679581782
transform 1 0 25248 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_264
timestamp 1679581782
transform 1 0 25920 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_271
timestamp 1679581782
transform 1 0 26592 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_278
timestamp 1679581782
transform 1 0 27264 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_285
timestamp 1679581782
transform 1 0 27936 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_292
timestamp 1679581782
transform 1 0 28608 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_299
timestamp 1679581782
transform 1 0 29280 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_306
timestamp 1679581782
transform 1 0 29952 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_313
timestamp 1679581782
transform 1 0 30624 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_320
timestamp 1679581782
transform 1 0 31296 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_327
timestamp 1679581782
transform 1 0 31968 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_334
timestamp 1679581782
transform 1 0 32640 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_341
timestamp 1679581782
transform 1 0 33312 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_348
timestamp 1679581782
transform 1 0 33984 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_355
timestamp 1679581782
transform 1 0 34656 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_362
timestamp 1679581782
transform 1 0 35328 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_369
timestamp 1679581782
transform 1 0 36000 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_376
timestamp 1679581782
transform 1 0 36672 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_383
timestamp 1679581782
transform 1 0 37344 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_390
timestamp 1679581782
transform 1 0 38016 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_397
timestamp 1679581782
transform 1 0 38688 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_404
timestamp 1679581782
transform 1 0 39360 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_411
timestamp 1679581782
transform 1 0 40032 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_418
timestamp 1679581782
transform 1 0 40704 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_425
timestamp 1679581782
transform 1 0 41376 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_432
timestamp 1679581782
transform 1 0 42048 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_439
timestamp 1679581782
transform 1 0 42720 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_446
timestamp 1679581782
transform 1 0 43392 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_453
timestamp 1679581782
transform 1 0 44064 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_460
timestamp 1679581782
transform 1 0 44736 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_467
timestamp 1679581782
transform 1 0 45408 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_474
timestamp 1679581782
transform 1 0 46080 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_481
timestamp 1679581782
transform 1 0 46752 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_488
timestamp 1679581782
transform 1 0 47424 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_495
timestamp 1679581782
transform 1 0 48096 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_502
timestamp 1679581782
transform 1 0 48768 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_509
timestamp 1679581782
transform 1 0 49440 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_516
timestamp 1679581782
transform 1 0 50112 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_523
timestamp 1679581782
transform 1 0 50784 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_530
timestamp 1679581782
transform 1 0 51456 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_537
timestamp 1679581782
transform 1 0 52128 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_544
timestamp 1679581782
transform 1 0 52800 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_551
timestamp 1679581782
transform 1 0 53472 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_558
timestamp 1679581782
transform 1 0 54144 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_565
timestamp 1679581782
transform 1 0 54816 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_572
timestamp 1679581782
transform 1 0 55488 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_579
timestamp 1679581782
transform 1 0 56160 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_586
timestamp 1679581782
transform 1 0 56832 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_593
timestamp 1679581782
transform 1 0 57504 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_600
timestamp 1679581782
transform 1 0 58176 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_607
timestamp 1679581782
transform 1 0 58848 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_614
timestamp 1679581782
transform 1 0 59520 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_621
timestamp 1679581782
transform 1 0 60192 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_628
timestamp 1679581782
transform 1 0 60864 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_635
timestamp 1679581782
transform 1 0 61536 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_642
timestamp 1679581782
transform 1 0 62208 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_649
timestamp 1679581782
transform 1 0 62880 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_656
timestamp 1679581782
transform 1 0 63552 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_663
timestamp 1679581782
transform 1 0 64224 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_670
timestamp 1679581782
transform 1 0 64896 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_677
timestamp 1679581782
transform 1 0 65568 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_684
timestamp 1679581782
transform 1 0 66240 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_691
timestamp 1679581782
transform 1 0 66912 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_698
timestamp 1679581782
transform 1 0 67584 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_705
timestamp 1679581782
transform 1 0 68256 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_712
timestamp 1679581782
transform 1 0 68928 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_719
timestamp 1679581782
transform 1 0 69600 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_726
timestamp 1679581782
transform 1 0 70272 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_733
timestamp 1679581782
transform 1 0 70944 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_740
timestamp 1679581782
transform 1 0 71616 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_747
timestamp 1679581782
transform 1 0 72288 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_754
timestamp 1679581782
transform 1 0 72960 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_761
timestamp 1679581782
transform 1 0 73632 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_768
timestamp 1679581782
transform 1 0 74304 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_775
timestamp 1679581782
transform 1 0 74976 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_782
timestamp 1679581782
transform 1 0 75648 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_789
timestamp 1679581782
transform 1 0 76320 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_796
timestamp 1679581782
transform 1 0 76992 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_803
timestamp 1679581782
transform 1 0 77664 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_810
timestamp 1679581782
transform 1 0 78336 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_817
timestamp 1679581782
transform 1 0 79008 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_824
timestamp 1679581782
transform 1 0 79680 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_831
timestamp 1679581782
transform 1 0 80352 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_838
timestamp 1679581782
transform 1 0 81024 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_845
timestamp 1679581782
transform 1 0 81696 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_852
timestamp 1679581782
transform 1 0 82368 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_859
timestamp 1679581782
transform 1 0 83040 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_866
timestamp 1679581782
transform 1 0 83712 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_873
timestamp 1679581782
transform 1 0 84384 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_880
timestamp 1679581782
transform 1 0 85056 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_887
timestamp 1679581782
transform 1 0 85728 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_894
timestamp 1679581782
transform 1 0 86400 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_901
timestamp 1679581782
transform 1 0 87072 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_908
timestamp 1679581782
transform 1 0 87744 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_915
timestamp 1679581782
transform 1 0 88416 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_922
timestamp 1679581782
transform 1 0 89088 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_929
timestamp 1679581782
transform 1 0 89760 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_936
timestamp 1679581782
transform 1 0 90432 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_943
timestamp 1679581782
transform 1 0 91104 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_950
timestamp 1679581782
transform 1 0 91776 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_957
timestamp 1679581782
transform 1 0 92448 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_964
timestamp 1679581782
transform 1 0 93120 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_971
timestamp 1679581782
transform 1 0 93792 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_978
timestamp 1679581782
transform 1 0 94464 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_985
timestamp 1679581782
transform 1 0 95136 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_992
timestamp 1679581782
transform 1 0 95808 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_999
timestamp 1679581782
transform 1 0 96480 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_1006
timestamp 1679581782
transform 1 0 97152 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_1013
timestamp 1679581782
transform 1 0 97824 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_1020
timestamp 1679581782
transform 1 0 98496 0 -1 35532
box -48 -56 720 834
use sg13g2_fill_2  FILLER_45_1027
timestamp 1677580104
transform 1 0 99168 0 -1 35532
box -48 -56 240 834
use sg13g2_decap_8  FILLER_46_0
timestamp 1679581782
transform 1 0 576 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_7
timestamp 1679581782
transform 1 0 1248 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_14
timestamp 1679581782
transform 1 0 1920 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_21
timestamp 1679581782
transform 1 0 2592 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_28
timestamp 1679581782
transform 1 0 3264 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_35
timestamp 1679581782
transform 1 0 3936 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_42
timestamp 1679581782
transform 1 0 4608 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_49
timestamp 1679581782
transform 1 0 5280 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_56
timestamp 1679581782
transform 1 0 5952 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_63
timestamp 1679581782
transform 1 0 6624 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_70
timestamp 1679581782
transform 1 0 7296 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_77
timestamp 1679581782
transform 1 0 7968 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_84
timestamp 1679581782
transform 1 0 8640 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_91
timestamp 1679581782
transform 1 0 9312 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_98
timestamp 1679581782
transform 1 0 9984 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_105
timestamp 1679581782
transform 1 0 10656 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_112
timestamp 1679581782
transform 1 0 11328 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_119
timestamp 1679581782
transform 1 0 12000 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_126
timestamp 1679581782
transform 1 0 12672 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_133
timestamp 1679581782
transform 1 0 13344 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_140
timestamp 1679581782
transform 1 0 14016 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_147
timestamp 1679581782
transform 1 0 14688 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_154
timestamp 1679581782
transform 1 0 15360 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_161
timestamp 1679581782
transform 1 0 16032 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_168
timestamp 1679581782
transform 1 0 16704 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_175
timestamp 1679581782
transform 1 0 17376 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_182
timestamp 1679581782
transform 1 0 18048 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_189
timestamp 1679581782
transform 1 0 18720 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_196
timestamp 1679581782
transform 1 0 19392 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_203
timestamp 1679581782
transform 1 0 20064 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_210
timestamp 1679581782
transform 1 0 20736 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_217
timestamp 1679581782
transform 1 0 21408 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_224
timestamp 1679581782
transform 1 0 22080 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_231
timestamp 1679581782
transform 1 0 22752 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_238
timestamp 1679581782
transform 1 0 23424 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_245
timestamp 1679581782
transform 1 0 24096 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_252
timestamp 1679581782
transform 1 0 24768 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_259
timestamp 1679581782
transform 1 0 25440 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_266
timestamp 1679581782
transform 1 0 26112 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_273
timestamp 1679581782
transform 1 0 26784 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_280
timestamp 1679581782
transform 1 0 27456 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_287
timestamp 1679581782
transform 1 0 28128 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_294
timestamp 1679581782
transform 1 0 28800 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_301
timestamp 1679581782
transform 1 0 29472 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_308
timestamp 1679581782
transform 1 0 30144 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_315
timestamp 1679581782
transform 1 0 30816 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_322
timestamp 1679581782
transform 1 0 31488 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_329
timestamp 1679581782
transform 1 0 32160 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_336
timestamp 1679581782
transform 1 0 32832 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_343
timestamp 1679581782
transform 1 0 33504 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_350
timestamp 1679581782
transform 1 0 34176 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_357
timestamp 1679581782
transform 1 0 34848 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_364
timestamp 1679581782
transform 1 0 35520 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_371
timestamp 1679581782
transform 1 0 36192 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_378
timestamp 1679581782
transform 1 0 36864 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_385
timestamp 1679581782
transform 1 0 37536 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_392
timestamp 1679581782
transform 1 0 38208 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_399
timestamp 1679581782
transform 1 0 38880 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_406
timestamp 1679581782
transform 1 0 39552 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_413
timestamp 1679581782
transform 1 0 40224 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_420
timestamp 1679581782
transform 1 0 40896 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_427
timestamp 1679581782
transform 1 0 41568 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_434
timestamp 1679581782
transform 1 0 42240 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_441
timestamp 1679581782
transform 1 0 42912 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_448
timestamp 1679581782
transform 1 0 43584 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_455
timestamp 1679581782
transform 1 0 44256 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_462
timestamp 1679581782
transform 1 0 44928 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_469
timestamp 1679581782
transform 1 0 45600 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_476
timestamp 1679581782
transform 1 0 46272 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_483
timestamp 1679581782
transform 1 0 46944 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_490
timestamp 1679581782
transform 1 0 47616 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_497
timestamp 1679581782
transform 1 0 48288 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_504
timestamp 1679581782
transform 1 0 48960 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_511
timestamp 1679581782
transform 1 0 49632 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_518
timestamp 1679581782
transform 1 0 50304 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_525
timestamp 1679581782
transform 1 0 50976 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_532
timestamp 1679581782
transform 1 0 51648 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_539
timestamp 1679581782
transform 1 0 52320 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_546
timestamp 1679581782
transform 1 0 52992 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_553
timestamp 1679581782
transform 1 0 53664 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_560
timestamp 1679581782
transform 1 0 54336 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_567
timestamp 1679581782
transform 1 0 55008 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_574
timestamp 1679581782
transform 1 0 55680 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_581
timestamp 1679581782
transform 1 0 56352 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_588
timestamp 1679581782
transform 1 0 57024 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_595
timestamp 1679581782
transform 1 0 57696 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_602
timestamp 1679581782
transform 1 0 58368 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_609
timestamp 1679581782
transform 1 0 59040 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_616
timestamp 1679581782
transform 1 0 59712 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_623
timestamp 1679581782
transform 1 0 60384 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_630
timestamp 1679581782
transform 1 0 61056 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_637
timestamp 1679581782
transform 1 0 61728 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_644
timestamp 1679581782
transform 1 0 62400 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_651
timestamp 1679581782
transform 1 0 63072 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_658
timestamp 1679581782
transform 1 0 63744 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_665
timestamp 1679581782
transform 1 0 64416 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_672
timestamp 1679581782
transform 1 0 65088 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_679
timestamp 1679581782
transform 1 0 65760 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_686
timestamp 1679581782
transform 1 0 66432 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_693
timestamp 1679581782
transform 1 0 67104 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_700
timestamp 1679581782
transform 1 0 67776 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_707
timestamp 1679581782
transform 1 0 68448 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_714
timestamp 1679581782
transform 1 0 69120 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_721
timestamp 1679581782
transform 1 0 69792 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_728
timestamp 1679581782
transform 1 0 70464 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_735
timestamp 1679581782
transform 1 0 71136 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_742
timestamp 1679581782
transform 1 0 71808 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_749
timestamp 1679581782
transform 1 0 72480 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_756
timestamp 1679581782
transform 1 0 73152 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_763
timestamp 1679581782
transform 1 0 73824 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_770
timestamp 1679581782
transform 1 0 74496 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_777
timestamp 1679581782
transform 1 0 75168 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_784
timestamp 1679581782
transform 1 0 75840 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_791
timestamp 1679581782
transform 1 0 76512 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_798
timestamp 1679581782
transform 1 0 77184 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_805
timestamp 1679581782
transform 1 0 77856 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_812
timestamp 1679581782
transform 1 0 78528 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_819
timestamp 1679581782
transform 1 0 79200 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_826
timestamp 1679581782
transform 1 0 79872 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_833
timestamp 1679581782
transform 1 0 80544 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_840
timestamp 1679581782
transform 1 0 81216 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_847
timestamp 1679581782
transform 1 0 81888 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_854
timestamp 1679581782
transform 1 0 82560 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_861
timestamp 1679581782
transform 1 0 83232 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_868
timestamp 1679581782
transform 1 0 83904 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_875
timestamp 1679581782
transform 1 0 84576 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_882
timestamp 1679581782
transform 1 0 85248 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_889
timestamp 1679581782
transform 1 0 85920 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_896
timestamp 1679581782
transform 1 0 86592 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_903
timestamp 1679581782
transform 1 0 87264 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_910
timestamp 1679581782
transform 1 0 87936 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_917
timestamp 1679581782
transform 1 0 88608 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_924
timestamp 1679581782
transform 1 0 89280 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_931
timestamp 1679581782
transform 1 0 89952 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_938
timestamp 1679581782
transform 1 0 90624 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_945
timestamp 1679581782
transform 1 0 91296 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_952
timestamp 1679581782
transform 1 0 91968 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_959
timestamp 1679581782
transform 1 0 92640 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_966
timestamp 1679581782
transform 1 0 93312 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_973
timestamp 1679581782
transform 1 0 93984 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_980
timestamp 1679581782
transform 1 0 94656 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_987
timestamp 1679581782
transform 1 0 95328 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_994
timestamp 1679581782
transform 1 0 96000 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_1001
timestamp 1679581782
transform 1 0 96672 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_1008
timestamp 1679581782
transform 1 0 97344 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_1015
timestamp 1679581782
transform 1 0 98016 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_1022
timestamp 1679581782
transform 1 0 98688 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_0
timestamp 1679581782
transform 1 0 576 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_7
timestamp 1679581782
transform 1 0 1248 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_14
timestamp 1679581782
transform 1 0 1920 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_21
timestamp 1679581782
transform 1 0 2592 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_28
timestamp 1679581782
transform 1 0 3264 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_35
timestamp 1679581782
transform 1 0 3936 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_42
timestamp 1679581782
transform 1 0 4608 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_49
timestamp 1679581782
transform 1 0 5280 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_56
timestamp 1679581782
transform 1 0 5952 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_63
timestamp 1679581782
transform 1 0 6624 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_70
timestamp 1679581782
transform 1 0 7296 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_77
timestamp 1679581782
transform 1 0 7968 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_84
timestamp 1679581782
transform 1 0 8640 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_91
timestamp 1679581782
transform 1 0 9312 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_98
timestamp 1679581782
transform 1 0 9984 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_105
timestamp 1679581782
transform 1 0 10656 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_112
timestamp 1679581782
transform 1 0 11328 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_119
timestamp 1679581782
transform 1 0 12000 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_126
timestamp 1679581782
transform 1 0 12672 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_133
timestamp 1679581782
transform 1 0 13344 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_140
timestamp 1679581782
transform 1 0 14016 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_147
timestamp 1679581782
transform 1 0 14688 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_154
timestamp 1679581782
transform 1 0 15360 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_161
timestamp 1679581782
transform 1 0 16032 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_168
timestamp 1679581782
transform 1 0 16704 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_175
timestamp 1679581782
transform 1 0 17376 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_182
timestamp 1679581782
transform 1 0 18048 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_189
timestamp 1679581782
transform 1 0 18720 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_196
timestamp 1679581782
transform 1 0 19392 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_203
timestamp 1679581782
transform 1 0 20064 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_210
timestamp 1679581782
transform 1 0 20736 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_217
timestamp 1679581782
transform 1 0 21408 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_224
timestamp 1679581782
transform 1 0 22080 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_231
timestamp 1679581782
transform 1 0 22752 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_238
timestamp 1679581782
transform 1 0 23424 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_245
timestamp 1679581782
transform 1 0 24096 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_252
timestamp 1679581782
transform 1 0 24768 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_259
timestamp 1679581782
transform 1 0 25440 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_266
timestamp 1679581782
transform 1 0 26112 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_273
timestamp 1679581782
transform 1 0 26784 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_280
timestamp 1679581782
transform 1 0 27456 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_287
timestamp 1679581782
transform 1 0 28128 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_294
timestamp 1679581782
transform 1 0 28800 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_301
timestamp 1679581782
transform 1 0 29472 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_308
timestamp 1679581782
transform 1 0 30144 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_315
timestamp 1679581782
transform 1 0 30816 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_322
timestamp 1679581782
transform 1 0 31488 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_329
timestamp 1679581782
transform 1 0 32160 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_336
timestamp 1679581782
transform 1 0 32832 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_343
timestamp 1679581782
transform 1 0 33504 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_350
timestamp 1679581782
transform 1 0 34176 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_357
timestamp 1679581782
transform 1 0 34848 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_364
timestamp 1679581782
transform 1 0 35520 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_371
timestamp 1679581782
transform 1 0 36192 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_378
timestamp 1679581782
transform 1 0 36864 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_385
timestamp 1679581782
transform 1 0 37536 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_392
timestamp 1679581782
transform 1 0 38208 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_399
timestamp 1679581782
transform 1 0 38880 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_406
timestamp 1679581782
transform 1 0 39552 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_413
timestamp 1679581782
transform 1 0 40224 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_420
timestamp 1679581782
transform 1 0 40896 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_427
timestamp 1679581782
transform 1 0 41568 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_434
timestamp 1679581782
transform 1 0 42240 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_441
timestamp 1679581782
transform 1 0 42912 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_448
timestamp 1679581782
transform 1 0 43584 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_455
timestamp 1679581782
transform 1 0 44256 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_462
timestamp 1679581782
transform 1 0 44928 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_469
timestamp 1679581782
transform 1 0 45600 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_476
timestamp 1679581782
transform 1 0 46272 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_483
timestamp 1679581782
transform 1 0 46944 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_490
timestamp 1679581782
transform 1 0 47616 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_497
timestamp 1679581782
transform 1 0 48288 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_504
timestamp 1679581782
transform 1 0 48960 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_511
timestamp 1679581782
transform 1 0 49632 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_518
timestamp 1679581782
transform 1 0 50304 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_525
timestamp 1679581782
transform 1 0 50976 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_532
timestamp 1679581782
transform 1 0 51648 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_539
timestamp 1679581782
transform 1 0 52320 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_546
timestamp 1679581782
transform 1 0 52992 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_553
timestamp 1679581782
transform 1 0 53664 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_560
timestamp 1679581782
transform 1 0 54336 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_567
timestamp 1679581782
transform 1 0 55008 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_574
timestamp 1679581782
transform 1 0 55680 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_581
timestamp 1679581782
transform 1 0 56352 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_588
timestamp 1679581782
transform 1 0 57024 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_595
timestamp 1679581782
transform 1 0 57696 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_602
timestamp 1679581782
transform 1 0 58368 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_609
timestamp 1679581782
transform 1 0 59040 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_616
timestamp 1679581782
transform 1 0 59712 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_623
timestamp 1679581782
transform 1 0 60384 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_630
timestamp 1679581782
transform 1 0 61056 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_637
timestamp 1679581782
transform 1 0 61728 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_644
timestamp 1679581782
transform 1 0 62400 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_651
timestamp 1679581782
transform 1 0 63072 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_658
timestamp 1679581782
transform 1 0 63744 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_665
timestamp 1679581782
transform 1 0 64416 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_672
timestamp 1679581782
transform 1 0 65088 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_679
timestamp 1679581782
transform 1 0 65760 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_686
timestamp 1679581782
transform 1 0 66432 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_693
timestamp 1679581782
transform 1 0 67104 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_700
timestamp 1679581782
transform 1 0 67776 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_707
timestamp 1679581782
transform 1 0 68448 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_714
timestamp 1679581782
transform 1 0 69120 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_721
timestamp 1679581782
transform 1 0 69792 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_728
timestamp 1679581782
transform 1 0 70464 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_735
timestamp 1679581782
transform 1 0 71136 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_742
timestamp 1679581782
transform 1 0 71808 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_749
timestamp 1679581782
transform 1 0 72480 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_756
timestamp 1679581782
transform 1 0 73152 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_763
timestamp 1679581782
transform 1 0 73824 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_770
timestamp 1679581782
transform 1 0 74496 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_777
timestamp 1679581782
transform 1 0 75168 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_784
timestamp 1679581782
transform 1 0 75840 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_791
timestamp 1679581782
transform 1 0 76512 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_798
timestamp 1679581782
transform 1 0 77184 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_805
timestamp 1679581782
transform 1 0 77856 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_812
timestamp 1679581782
transform 1 0 78528 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_819
timestamp 1679581782
transform 1 0 79200 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_826
timestamp 1679581782
transform 1 0 79872 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_833
timestamp 1679581782
transform 1 0 80544 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_840
timestamp 1679581782
transform 1 0 81216 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_847
timestamp 1679581782
transform 1 0 81888 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_854
timestamp 1679581782
transform 1 0 82560 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_861
timestamp 1679581782
transform 1 0 83232 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_868
timestamp 1679581782
transform 1 0 83904 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_875
timestamp 1679581782
transform 1 0 84576 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_882
timestamp 1679581782
transform 1 0 85248 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_889
timestamp 1679581782
transform 1 0 85920 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_896
timestamp 1679581782
transform 1 0 86592 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_903
timestamp 1679581782
transform 1 0 87264 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_910
timestamp 1679581782
transform 1 0 87936 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_917
timestamp 1679581782
transform 1 0 88608 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_924
timestamp 1679581782
transform 1 0 89280 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_931
timestamp 1679581782
transform 1 0 89952 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_938
timestamp 1679581782
transform 1 0 90624 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_945
timestamp 1679581782
transform 1 0 91296 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_952
timestamp 1679581782
transform 1 0 91968 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_959
timestamp 1679581782
transform 1 0 92640 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_966
timestamp 1679581782
transform 1 0 93312 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_973
timestamp 1679581782
transform 1 0 93984 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_980
timestamp 1679581782
transform 1 0 94656 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_987
timestamp 1679581782
transform 1 0 95328 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_994
timestamp 1679581782
transform 1 0 96000 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_1001
timestamp 1679581782
transform 1 0 96672 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_1008
timestamp 1679581782
transform 1 0 97344 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_1015
timestamp 1679581782
transform 1 0 98016 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_1022
timestamp 1679581782
transform 1 0 98688 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_0
timestamp 1679581782
transform 1 0 576 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_7
timestamp 1679581782
transform 1 0 1248 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_14
timestamp 1679581782
transform 1 0 1920 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_21
timestamp 1679581782
transform 1 0 2592 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_28
timestamp 1679581782
transform 1 0 3264 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_35
timestamp 1679581782
transform 1 0 3936 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_42
timestamp 1679581782
transform 1 0 4608 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_49
timestamp 1679581782
transform 1 0 5280 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_56
timestamp 1679581782
transform 1 0 5952 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_63
timestamp 1679581782
transform 1 0 6624 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_70
timestamp 1679581782
transform 1 0 7296 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_77
timestamp 1679581782
transform 1 0 7968 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_84
timestamp 1679581782
transform 1 0 8640 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_91
timestamp 1679581782
transform 1 0 9312 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_98
timestamp 1679581782
transform 1 0 9984 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_105
timestamp 1679581782
transform 1 0 10656 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_112
timestamp 1679581782
transform 1 0 11328 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_119
timestamp 1679581782
transform 1 0 12000 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_126
timestamp 1679581782
transform 1 0 12672 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_133
timestamp 1679581782
transform 1 0 13344 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_140
timestamp 1679581782
transform 1 0 14016 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_147
timestamp 1679581782
transform 1 0 14688 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_154
timestamp 1679581782
transform 1 0 15360 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_161
timestamp 1679581782
transform 1 0 16032 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_168
timestamp 1679581782
transform 1 0 16704 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_175
timestamp 1679581782
transform 1 0 17376 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_182
timestamp 1679581782
transform 1 0 18048 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_189
timestamp 1679581782
transform 1 0 18720 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_196
timestamp 1679581782
transform 1 0 19392 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_203
timestamp 1679581782
transform 1 0 20064 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_210
timestamp 1679581782
transform 1 0 20736 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_217
timestamp 1679581782
transform 1 0 21408 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_224
timestamp 1679581782
transform 1 0 22080 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_231
timestamp 1679581782
transform 1 0 22752 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_238
timestamp 1679581782
transform 1 0 23424 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_245
timestamp 1679581782
transform 1 0 24096 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_252
timestamp 1679581782
transform 1 0 24768 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_259
timestamp 1679581782
transform 1 0 25440 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_266
timestamp 1679581782
transform 1 0 26112 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_273
timestamp 1679581782
transform 1 0 26784 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_280
timestamp 1679581782
transform 1 0 27456 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_287
timestamp 1679581782
transform 1 0 28128 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_294
timestamp 1679581782
transform 1 0 28800 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_301
timestamp 1679581782
transform 1 0 29472 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_308
timestamp 1679581782
transform 1 0 30144 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_315
timestamp 1679581782
transform 1 0 30816 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_322
timestamp 1679581782
transform 1 0 31488 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_329
timestamp 1679581782
transform 1 0 32160 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_336
timestamp 1679581782
transform 1 0 32832 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_343
timestamp 1679581782
transform 1 0 33504 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_350
timestamp 1679581782
transform 1 0 34176 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_357
timestamp 1679581782
transform 1 0 34848 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_364
timestamp 1679581782
transform 1 0 35520 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_371
timestamp 1679581782
transform 1 0 36192 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_378
timestamp 1679581782
transform 1 0 36864 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_385
timestamp 1679581782
transform 1 0 37536 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_392
timestamp 1679581782
transform 1 0 38208 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_399
timestamp 1679581782
transform 1 0 38880 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_406
timestamp 1679581782
transform 1 0 39552 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_413
timestamp 1679581782
transform 1 0 40224 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_420
timestamp 1679581782
transform 1 0 40896 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_427
timestamp 1679581782
transform 1 0 41568 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_434
timestamp 1679581782
transform 1 0 42240 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_441
timestamp 1679581782
transform 1 0 42912 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_448
timestamp 1679581782
transform 1 0 43584 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_455
timestamp 1679581782
transform 1 0 44256 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_462
timestamp 1679581782
transform 1 0 44928 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_469
timestamp 1679581782
transform 1 0 45600 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_476
timestamp 1679581782
transform 1 0 46272 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_483
timestamp 1679581782
transform 1 0 46944 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_490
timestamp 1679581782
transform 1 0 47616 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_497
timestamp 1679581782
transform 1 0 48288 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_504
timestamp 1679581782
transform 1 0 48960 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_511
timestamp 1679581782
transform 1 0 49632 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_518
timestamp 1679581782
transform 1 0 50304 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_525
timestamp 1679581782
transform 1 0 50976 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_532
timestamp 1679581782
transform 1 0 51648 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_539
timestamp 1679581782
transform 1 0 52320 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_546
timestamp 1679581782
transform 1 0 52992 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_553
timestamp 1679581782
transform 1 0 53664 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_560
timestamp 1679581782
transform 1 0 54336 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_567
timestamp 1679581782
transform 1 0 55008 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_574
timestamp 1679581782
transform 1 0 55680 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_581
timestamp 1679581782
transform 1 0 56352 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_588
timestamp 1679581782
transform 1 0 57024 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_595
timestamp 1679581782
transform 1 0 57696 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_602
timestamp 1679581782
transform 1 0 58368 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_609
timestamp 1679581782
transform 1 0 59040 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_616
timestamp 1679581782
transform 1 0 59712 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_623
timestamp 1679581782
transform 1 0 60384 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_630
timestamp 1679581782
transform 1 0 61056 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_637
timestamp 1679581782
transform 1 0 61728 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_644
timestamp 1679581782
transform 1 0 62400 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_651
timestamp 1679581782
transform 1 0 63072 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_658
timestamp 1679581782
transform 1 0 63744 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_665
timestamp 1679581782
transform 1 0 64416 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_672
timestamp 1679581782
transform 1 0 65088 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_679
timestamp 1679581782
transform 1 0 65760 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_686
timestamp 1679581782
transform 1 0 66432 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_693
timestamp 1679581782
transform 1 0 67104 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_700
timestamp 1679581782
transform 1 0 67776 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_707
timestamp 1679581782
transform 1 0 68448 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_714
timestamp 1679581782
transform 1 0 69120 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_721
timestamp 1679581782
transform 1 0 69792 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_728
timestamp 1679581782
transform 1 0 70464 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_735
timestamp 1679581782
transform 1 0 71136 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_742
timestamp 1679581782
transform 1 0 71808 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_749
timestamp 1679581782
transform 1 0 72480 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_756
timestamp 1679581782
transform 1 0 73152 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_763
timestamp 1679581782
transform 1 0 73824 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_770
timestamp 1679581782
transform 1 0 74496 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_777
timestamp 1679581782
transform 1 0 75168 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_784
timestamp 1679581782
transform 1 0 75840 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_791
timestamp 1679581782
transform 1 0 76512 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_798
timestamp 1679581782
transform 1 0 77184 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_805
timestamp 1679581782
transform 1 0 77856 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_812
timestamp 1679581782
transform 1 0 78528 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_819
timestamp 1679581782
transform 1 0 79200 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_826
timestamp 1679581782
transform 1 0 79872 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_833
timestamp 1679581782
transform 1 0 80544 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_840
timestamp 1679581782
transform 1 0 81216 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_847
timestamp 1679581782
transform 1 0 81888 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_854
timestamp 1679581782
transform 1 0 82560 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_861
timestamp 1679581782
transform 1 0 83232 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_868
timestamp 1679581782
transform 1 0 83904 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_875
timestamp 1679581782
transform 1 0 84576 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_882
timestamp 1679581782
transform 1 0 85248 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_889
timestamp 1679581782
transform 1 0 85920 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_896
timestamp 1679581782
transform 1 0 86592 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_903
timestamp 1679581782
transform 1 0 87264 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_910
timestamp 1679581782
transform 1 0 87936 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_917
timestamp 1679581782
transform 1 0 88608 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_924
timestamp 1679581782
transform 1 0 89280 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_931
timestamp 1679581782
transform 1 0 89952 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_938
timestamp 1679581782
transform 1 0 90624 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_945
timestamp 1679581782
transform 1 0 91296 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_952
timestamp 1679581782
transform 1 0 91968 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_959
timestamp 1679581782
transform 1 0 92640 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_966
timestamp 1679581782
transform 1 0 93312 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_973
timestamp 1679581782
transform 1 0 93984 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_980
timestamp 1679581782
transform 1 0 94656 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_987
timestamp 1679581782
transform 1 0 95328 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_994
timestamp 1679581782
transform 1 0 96000 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_1001
timestamp 1679581782
transform 1 0 96672 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_1008
timestamp 1679581782
transform 1 0 97344 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_1015
timestamp 1679581782
transform 1 0 98016 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_1022
timestamp 1679581782
transform 1 0 98688 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_0
timestamp 1679581782
transform 1 0 576 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_7
timestamp 1679581782
transform 1 0 1248 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_14
timestamp 1679581782
transform 1 0 1920 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_21
timestamp 1679581782
transform 1 0 2592 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_28
timestamp 1679581782
transform 1 0 3264 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_35
timestamp 1679581782
transform 1 0 3936 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_42
timestamp 1679581782
transform 1 0 4608 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_49
timestamp 1679581782
transform 1 0 5280 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_56
timestamp 1679581782
transform 1 0 5952 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_63
timestamp 1679581782
transform 1 0 6624 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_70
timestamp 1679581782
transform 1 0 7296 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_77
timestamp 1679581782
transform 1 0 7968 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_84
timestamp 1679581782
transform 1 0 8640 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_91
timestamp 1679581782
transform 1 0 9312 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_98
timestamp 1679581782
transform 1 0 9984 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_105
timestamp 1679581782
transform 1 0 10656 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_112
timestamp 1679581782
transform 1 0 11328 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_119
timestamp 1679581782
transform 1 0 12000 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_126
timestamp 1679581782
transform 1 0 12672 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_133
timestamp 1679581782
transform 1 0 13344 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_140
timestamp 1679581782
transform 1 0 14016 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_147
timestamp 1679581782
transform 1 0 14688 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_154
timestamp 1679581782
transform 1 0 15360 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_161
timestamp 1679581782
transform 1 0 16032 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_168
timestamp 1679581782
transform 1 0 16704 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_175
timestamp 1679581782
transform 1 0 17376 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_182
timestamp 1679581782
transform 1 0 18048 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_189
timestamp 1679581782
transform 1 0 18720 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_196
timestamp 1679581782
transform 1 0 19392 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_203
timestamp 1679581782
transform 1 0 20064 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_210
timestamp 1679581782
transform 1 0 20736 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_217
timestamp 1679581782
transform 1 0 21408 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_224
timestamp 1679581782
transform 1 0 22080 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_231
timestamp 1679581782
transform 1 0 22752 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_238
timestamp 1679581782
transform 1 0 23424 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_245
timestamp 1679581782
transform 1 0 24096 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_252
timestamp 1679581782
transform 1 0 24768 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_259
timestamp 1679581782
transform 1 0 25440 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_266
timestamp 1679581782
transform 1 0 26112 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_273
timestamp 1679581782
transform 1 0 26784 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_280
timestamp 1679581782
transform 1 0 27456 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_287
timestamp 1679581782
transform 1 0 28128 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_294
timestamp 1679581782
transform 1 0 28800 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_301
timestamp 1679581782
transform 1 0 29472 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_308
timestamp 1679581782
transform 1 0 30144 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_315
timestamp 1679581782
transform 1 0 30816 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_322
timestamp 1679581782
transform 1 0 31488 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_329
timestamp 1679581782
transform 1 0 32160 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_336
timestamp 1679581782
transform 1 0 32832 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_343
timestamp 1679581782
transform 1 0 33504 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_350
timestamp 1679581782
transform 1 0 34176 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_357
timestamp 1679581782
transform 1 0 34848 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_364
timestamp 1679581782
transform 1 0 35520 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_371
timestamp 1679581782
transform 1 0 36192 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_378
timestamp 1679581782
transform 1 0 36864 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_385
timestamp 1679581782
transform 1 0 37536 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_392
timestamp 1679581782
transform 1 0 38208 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_399
timestamp 1679581782
transform 1 0 38880 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_406
timestamp 1679581782
transform 1 0 39552 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_413
timestamp 1679581782
transform 1 0 40224 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_420
timestamp 1679581782
transform 1 0 40896 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_427
timestamp 1679581782
transform 1 0 41568 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_434
timestamp 1679581782
transform 1 0 42240 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_441
timestamp 1679581782
transform 1 0 42912 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_448
timestamp 1679581782
transform 1 0 43584 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_455
timestamp 1679581782
transform 1 0 44256 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_462
timestamp 1679581782
transform 1 0 44928 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_469
timestamp 1679581782
transform 1 0 45600 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_476
timestamp 1679581782
transform 1 0 46272 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_483
timestamp 1679581782
transform 1 0 46944 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_490
timestamp 1679581782
transform 1 0 47616 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_497
timestamp 1679581782
transform 1 0 48288 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_504
timestamp 1679581782
transform 1 0 48960 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_511
timestamp 1679581782
transform 1 0 49632 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_518
timestamp 1679581782
transform 1 0 50304 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_525
timestamp 1679581782
transform 1 0 50976 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_532
timestamp 1679581782
transform 1 0 51648 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_539
timestamp 1679581782
transform 1 0 52320 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_546
timestamp 1679581782
transform 1 0 52992 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_553
timestamp 1679581782
transform 1 0 53664 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_560
timestamp 1679581782
transform 1 0 54336 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_567
timestamp 1679581782
transform 1 0 55008 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_574
timestamp 1679581782
transform 1 0 55680 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_581
timestamp 1679581782
transform 1 0 56352 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_588
timestamp 1679581782
transform 1 0 57024 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_595
timestamp 1679581782
transform 1 0 57696 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_602
timestamp 1679581782
transform 1 0 58368 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_609
timestamp 1679581782
transform 1 0 59040 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_616
timestamp 1679581782
transform 1 0 59712 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_623
timestamp 1679581782
transform 1 0 60384 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_630
timestamp 1679581782
transform 1 0 61056 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_637
timestamp 1679581782
transform 1 0 61728 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_644
timestamp 1679581782
transform 1 0 62400 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_651
timestamp 1679581782
transform 1 0 63072 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_658
timestamp 1679581782
transform 1 0 63744 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_665
timestamp 1679581782
transform 1 0 64416 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_672
timestamp 1679581782
transform 1 0 65088 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_679
timestamp 1679581782
transform 1 0 65760 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_686
timestamp 1679581782
transform 1 0 66432 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_693
timestamp 1679581782
transform 1 0 67104 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_700
timestamp 1679581782
transform 1 0 67776 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_707
timestamp 1679581782
transform 1 0 68448 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_714
timestamp 1679581782
transform 1 0 69120 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_721
timestamp 1679581782
transform 1 0 69792 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_728
timestamp 1679581782
transform 1 0 70464 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_735
timestamp 1679581782
transform 1 0 71136 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_742
timestamp 1679581782
transform 1 0 71808 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_749
timestamp 1679581782
transform 1 0 72480 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_756
timestamp 1679581782
transform 1 0 73152 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_763
timestamp 1679581782
transform 1 0 73824 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_770
timestamp 1679581782
transform 1 0 74496 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_777
timestamp 1679581782
transform 1 0 75168 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_784
timestamp 1679581782
transform 1 0 75840 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_791
timestamp 1679581782
transform 1 0 76512 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_798
timestamp 1679581782
transform 1 0 77184 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_805
timestamp 1679581782
transform 1 0 77856 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_812
timestamp 1679581782
transform 1 0 78528 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_819
timestamp 1679581782
transform 1 0 79200 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_826
timestamp 1679581782
transform 1 0 79872 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_833
timestamp 1679581782
transform 1 0 80544 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_840
timestamp 1679581782
transform 1 0 81216 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_847
timestamp 1679581782
transform 1 0 81888 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_854
timestamp 1679581782
transform 1 0 82560 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_861
timestamp 1679581782
transform 1 0 83232 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_868
timestamp 1679581782
transform 1 0 83904 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_875
timestamp 1679581782
transform 1 0 84576 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_882
timestamp 1679581782
transform 1 0 85248 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_889
timestamp 1679581782
transform 1 0 85920 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_896
timestamp 1679581782
transform 1 0 86592 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_903
timestamp 1679581782
transform 1 0 87264 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_910
timestamp 1679581782
transform 1 0 87936 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_917
timestamp 1679581782
transform 1 0 88608 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_924
timestamp 1679581782
transform 1 0 89280 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_931
timestamp 1679581782
transform 1 0 89952 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_938
timestamp 1679581782
transform 1 0 90624 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_945
timestamp 1679581782
transform 1 0 91296 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_952
timestamp 1679581782
transform 1 0 91968 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_959
timestamp 1679581782
transform 1 0 92640 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_966
timestamp 1679581782
transform 1 0 93312 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_973
timestamp 1679581782
transform 1 0 93984 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_980
timestamp 1679581782
transform 1 0 94656 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_987
timestamp 1679581782
transform 1 0 95328 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_994
timestamp 1679581782
transform 1 0 96000 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_1001
timestamp 1679581782
transform 1 0 96672 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_1008
timestamp 1679581782
transform 1 0 97344 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_1015
timestamp 1679581782
transform 1 0 98016 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_1022
timestamp 1679581782
transform 1 0 98688 0 -1 38556
box -48 -56 720 834
use sg13g2_tielo  heichips25_template_28
timestamp 1680000637
transform -1 0 960 0 -1 12852
box -48 -56 432 834
use sg13g2_tielo  heichips25_template_29
timestamp 1680000637
transform -1 0 960 0 1 12852
box -48 -56 432 834
use sg13g2_tielo  heichips25_template_30
timestamp 1680000637
transform -1 0 960 0 1 14364
box -48 -56 432 834
use sg13g2_tielo  heichips25_template_31
timestamp 1680000637
transform -1 0 960 0 -1 15876
box -48 -56 432 834
use sg13g2_tiehi  heichips25_template_33
timestamp 1680000651
transform -1 0 960 0 1 15876
box -48 -56 432 834
use sg13g2_tiehi  heichips25_template_34
timestamp 1680000651
transform -1 0 960 0 -1 17388
box -48 -56 432 834
use sg13g2_tiehi  heichips25_template_35
timestamp 1680000651
transform -1 0 960 0 1 17388
box -48 -56 432 834
use sg13g2_tiehi  heichips25_template_36
timestamp 1680000651
transform -1 0 960 0 -1 18900
box -48 -56 432 834
use sg13g2_tiehi  heichips25_template_37
timestamp 1680000651
transform -1 0 960 0 1 18900
box -48 -56 432 834
use sg13g2_tiehi  heichips25_template_38
timestamp 1680000651
transform -1 0 960 0 -1 20412
box -48 -56 432 834
use sg13g2_tiehi  heichips25_template_39
timestamp 1680000651
transform -1 0 960 0 1 20412
box -48 -56 432 834
use sg13g2_tiehi  heichips25_template_40
timestamp 1680000651
transform -1 0 960 0 1 21924
box -48 -56 432 834
use sg13g2_dlygate4sd3_1  hold1
timestamp 1677672058
transform -1 0 39360 0 1 15876
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold2
timestamp 1677672058
transform -1 0 29184 0 -1 18900
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold3
timestamp 1677672058
transform -1 0 40032 0 -1 20412
box -48 -56 912 834
use sg13g2_buf_2  input1
timestamp 1676381867
transform -1 0 1056 0 1 23436
box -48 -56 528 834
use sg13g2_buf_2  input2
timestamp 1676381867
transform -1 0 1056 0 -1 24948
box -48 -56 528 834
use sg13g2_buf_2  input3
timestamp 1676381867
transform -1 0 1056 0 1 24948
box -48 -56 528 834
use sg13g2_buf_2  input4
timestamp 1676381867
transform -1 0 1056 0 -1 26460
box -48 -56 528 834
use sg13g2_buf_2  input5
timestamp 1676381867
transform -1 0 1056 0 1 26460
box -48 -56 528 834
use sg13g2_buf_2  input6
timestamp 1676381867
transform -1 0 1056 0 -1 27972
box -48 -56 528 834
use sg13g2_buf_2  input7
timestamp 1676381867
transform -1 0 1056 0 1 27972
box -48 -56 528 834
use sg13g2_buf_1  input8
timestamp 1676381911
transform 1 0 576 0 1 29484
box -48 -56 432 834
use sg13g2_buf_1  input9
timestamp 1676381911
transform 1 0 576 0 -1 30996
box -48 -56 432 834
use sg13g2_buf_1  input10
timestamp 1676381911
transform 1 0 576 0 1 30996
box -48 -56 432 834
use sg13g2_buf_1  input11
timestamp 1676381911
transform 1 0 576 0 -1 32508
box -48 -56 432 834
use sg13g2_buf_2  input12
timestamp 1676381867
transform -1 0 1056 0 1 32508
box -48 -56 528 834
use sg13g2_buf_2  input13
timestamp 1676381867
transform -1 0 1056 0 -1 34020
box -48 -56 528 834
use sg13g2_buf_2  input14
timestamp 1676381867
transform -1 0 1056 0 1 34020
box -48 -56 528 834
use sg13g2_buf_2  input15
timestamp 1676381867
transform -1 0 1056 0 -1 35532
box -48 -56 528 834
use sg13g2_buf_1  output16
timestamp 1676381911
transform -1 0 960 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  output17
timestamp 1676381911
transform -1 0 960 0 1 9828
box -48 -56 432 834
use sg13g2_buf_1  output18
timestamp 1676381911
transform -1 0 960 0 -1 11340
box -48 -56 432 834
use sg13g2_buf_1  output19
timestamp 1676381911
transform -1 0 960 0 1 11340
box -48 -56 432 834
use sg13g2_buf_1  output20
timestamp 1676381911
transform -1 0 960 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  output21
timestamp 1676381911
transform -1 0 960 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  output22
timestamp 1676381911
transform -1 0 960 0 1 3780
box -48 -56 432 834
use sg13g2_buf_1  output23
timestamp 1676381911
transform -1 0 960 0 -1 5292
box -48 -56 432 834
use sg13g2_buf_1  output24
timestamp 1676381911
transform -1 0 960 0 1 5292
box -48 -56 432 834
use sg13g2_buf_1  output25
timestamp 1676381911
transform -1 0 960 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  output26
timestamp 1676381911
transform -1 0 960 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  output27
timestamp 1676381911
transform -1 0 960 0 1 8316
box -48 -56 432 834
<< labels >>
flabel metal6 s 4316 630 4756 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 19436 630 19876 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 34556 630 34996 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 49676 630 50116 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 64796 630 65236 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 79916 630 80356 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 95036 630 95476 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 3076 712 3516 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 18196 712 18636 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 33316 712 33756 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 48436 712 48876 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 63556 712 63996 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 78676 712 79116 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 93796 712 94236 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 36668 80 36748 0 FreeSans 320 0 0 0 clk
port 2 nsew signal input
flabel metal3 s 0 35828 80 35908 0 FreeSans 320 0 0 0 ena
port 3 nsew signal input
flabel metal3 s 0 37508 80 37588 0 FreeSans 320 0 0 0 rst_n
port 4 nsew signal input
flabel metal3 s 0 22388 80 22468 0 FreeSans 320 0 0 0 ui_in[0]
port 5 nsew signal input
flabel metal3 s 0 23228 80 23308 0 FreeSans 320 0 0 0 ui_in[1]
port 6 nsew signal input
flabel metal3 s 0 24068 80 24148 0 FreeSans 320 0 0 0 ui_in[2]
port 7 nsew signal input
flabel metal3 s 0 24908 80 24988 0 FreeSans 320 0 0 0 ui_in[3]
port 8 nsew signal input
flabel metal3 s 0 25748 80 25828 0 FreeSans 320 0 0 0 ui_in[4]
port 9 nsew signal input
flabel metal3 s 0 26588 80 26668 0 FreeSans 320 0 0 0 ui_in[5]
port 10 nsew signal input
flabel metal3 s 0 27428 80 27508 0 FreeSans 320 0 0 0 ui_in[6]
port 11 nsew signal input
flabel metal3 s 0 28268 80 28348 0 FreeSans 320 0 0 0 ui_in[7]
port 12 nsew signal input
flabel metal3 s 0 29108 80 29188 0 FreeSans 320 0 0 0 uio_in[0]
port 13 nsew signal input
flabel metal3 s 0 29948 80 30028 0 FreeSans 320 0 0 0 uio_in[1]
port 14 nsew signal input
flabel metal3 s 0 30788 80 30868 0 FreeSans 320 0 0 0 uio_in[2]
port 15 nsew signal input
flabel metal3 s 0 31628 80 31708 0 FreeSans 320 0 0 0 uio_in[3]
port 16 nsew signal input
flabel metal3 s 0 32468 80 32548 0 FreeSans 320 0 0 0 uio_in[4]
port 17 nsew signal input
flabel metal3 s 0 33308 80 33388 0 FreeSans 320 0 0 0 uio_in[5]
port 18 nsew signal input
flabel metal3 s 0 34148 80 34228 0 FreeSans 320 0 0 0 uio_in[6]
port 19 nsew signal input
flabel metal3 s 0 34988 80 35068 0 FreeSans 320 0 0 0 uio_in[7]
port 20 nsew signal input
flabel metal3 s 0 15668 80 15748 0 FreeSans 320 0 0 0 uio_oe[0]
port 21 nsew signal output
flabel metal3 s 0 16508 80 16588 0 FreeSans 320 0 0 0 uio_oe[1]
port 22 nsew signal output
flabel metal3 s 0 17348 80 17428 0 FreeSans 320 0 0 0 uio_oe[2]
port 23 nsew signal output
flabel metal3 s 0 18188 80 18268 0 FreeSans 320 0 0 0 uio_oe[3]
port 24 nsew signal output
flabel metal3 s 0 19028 80 19108 0 FreeSans 320 0 0 0 uio_oe[4]
port 25 nsew signal output
flabel metal3 s 0 19868 80 19948 0 FreeSans 320 0 0 0 uio_oe[5]
port 26 nsew signal output
flabel metal3 s 0 20708 80 20788 0 FreeSans 320 0 0 0 uio_oe[6]
port 27 nsew signal output
flabel metal3 s 0 21548 80 21628 0 FreeSans 320 0 0 0 uio_oe[7]
port 28 nsew signal output
flabel metal3 s 0 8948 80 9028 0 FreeSans 320 0 0 0 uio_out[0]
port 29 nsew signal output
flabel metal3 s 0 9788 80 9868 0 FreeSans 320 0 0 0 uio_out[1]
port 30 nsew signal output
flabel metal3 s 0 10628 80 10708 0 FreeSans 320 0 0 0 uio_out[2]
port 31 nsew signal output
flabel metal3 s 0 11468 80 11548 0 FreeSans 320 0 0 0 uio_out[3]
port 32 nsew signal output
flabel metal3 s 0 12308 80 12388 0 FreeSans 320 0 0 0 uio_out[4]
port 33 nsew signal output
flabel metal3 s 0 13148 80 13228 0 FreeSans 320 0 0 0 uio_out[5]
port 34 nsew signal output
flabel metal3 s 0 13988 80 14068 0 FreeSans 320 0 0 0 uio_out[6]
port 35 nsew signal output
flabel metal3 s 0 14828 80 14908 0 FreeSans 320 0 0 0 uio_out[7]
port 36 nsew signal output
flabel metal3 s 0 2228 80 2308 0 FreeSans 320 0 0 0 uo_out[0]
port 37 nsew signal output
flabel metal3 s 0 3068 80 3148 0 FreeSans 320 0 0 0 uo_out[1]
port 38 nsew signal output
flabel metal3 s 0 3908 80 3988 0 FreeSans 320 0 0 0 uo_out[2]
port 39 nsew signal output
flabel metal3 s 0 4748 80 4828 0 FreeSans 320 0 0 0 uo_out[3]
port 40 nsew signal output
flabel metal3 s 0 5588 80 5668 0 FreeSans 320 0 0 0 uo_out[4]
port 41 nsew signal output
flabel metal3 s 0 6428 80 6508 0 FreeSans 320 0 0 0 uo_out[5]
port 42 nsew signal output
flabel metal3 s 0 7268 80 7348 0 FreeSans 320 0 0 0 uo_out[6]
port 43 nsew signal output
flabel metal3 s 0 8108 80 8188 0 FreeSans 320 0 0 0 uo_out[7]
port 44 nsew signal output
rlabel via1 49968 38556 49968 38556 0 VGND
rlabel metal1 49968 37800 49968 37800 0 VPWR
rlabel metal2 27360 30870 27360 30870 0 Demo1.epsk_de1.bit_out\[0\]
rlabel metal3 36624 27048 36624 27048 0 Demo1.epsk_de1.bit_out\[1\]
rlabel metal2 18432 27888 18432 27888 0 Demo1.epsk_de1.bit_out\[2\]
rlabel metal3 27216 30660 27216 30660 0 Demo1.qam16_bits\[0\]
rlabel metal2 35616 29778 35616 29778 0 Demo1.qam16_bits\[1\]
rlabel metal2 17280 26964 17280 26964 0 Demo1.qam16_bits\[2\]
rlabel metal2 33792 16296 33792 16296 0 Demo1.qam16_bits\[3\]
rlabel metal2 19200 22050 19200 22050 0 _000_
rlabel metal2 21408 29904 21408 29904 0 _001_
rlabel metal2 34944 27048 34944 27048 0 _002_
rlabel metal3 18912 28308 18912 28308 0 _003_
rlabel metal2 29184 30744 29184 30744 0 _004_
rlabel metal2 31296 29778 31296 29778 0 _005_
rlabel metal2 15456 15918 15456 15918 0 _006_
rlabel metal2 23424 21462 23424 21462 0 _007_
rlabel metal2 34080 21336 34080 21336 0 _008_
rlabel metal2 22944 17808 22944 17808 0 _009_
rlabel metal2 22512 16884 22512 16884 0 _010_
rlabel metal2 14880 26418 14880 26418 0 _011_
rlabel metal2 37056 15834 37056 15834 0 _012_
rlabel metal2 38784 19320 38784 19320 0 _013_
rlabel metal3 26544 17724 26544 17724 0 _014_
rlabel metal2 34272 17346 34272 17346 0 _015_
rlabel metal2 28080 12432 28080 12432 0 _016_
rlabel metal2 27840 12642 27840 12642 0 _017_
rlabel metal2 27264 12558 27264 12558 0 _018_
rlabel metal2 22848 17682 22848 17682 0 _019_
rlabel metal2 22080 20286 22080 20286 0 _020_
rlabel metal2 16032 17304 16032 17304 0 _021_
rlabel metal2 22848 20454 22848 20454 0 _022_
rlabel metal3 29664 28308 29664 28308 0 _023_
rlabel metal2 29952 27678 29952 27678 0 _024_
rlabel metal2 28512 28224 28512 28224 0 _025_
rlabel metal2 29472 27090 29472 27090 0 _026_
rlabel metal2 28224 28434 28224 28434 0 _027_
rlabel metal3 27504 27720 27504 27720 0 _028_
rlabel metal2 28128 26712 28128 26712 0 _029_
rlabel metal3 22848 27804 22848 27804 0 _030_
rlabel metal2 22560 27901 22560 27901 0 _031_
rlabel metal3 21840 17976 21840 17976 0 _032_
rlabel metal2 28608 22260 28608 22260 0 _033_
rlabel metal2 28896 22344 28896 22344 0 _034_
rlabel metal2 26112 18606 26112 18606 0 _035_
rlabel metal2 26400 25830 26400 25830 0 _036_
rlabel metal3 21216 26796 21216 26796 0 _037_
rlabel metal2 20544 27090 20544 27090 0 _038_
rlabel metal2 22656 19530 22656 19530 0 _039_
rlabel metal2 19392 19068 19392 19068 0 _040_
rlabel metal2 18384 15456 18384 15456 0 _041_
rlabel metal2 27456 31332 27456 31332 0 _042_
rlabel metal3 36144 28980 36144 28980 0 _043_
rlabel metal2 18720 27510 18720 27510 0 _044_
rlabel metal3 34320 20076 34320 20076 0 _045_
rlabel metal2 33984 16674 33984 16674 0 _046_
rlabel metal3 30144 20832 30144 20832 0 _047_
rlabel metal2 30816 20874 30816 20874 0 _048_
rlabel metal2 34752 22218 34752 22218 0 _049_
rlabel metal2 34840 22134 34840 22134 0 _050_
rlabel metal2 34176 22428 34176 22428 0 _051_
rlabel metal3 33312 22260 33312 22260 0 _052_
rlabel metal2 35040 22218 35040 22218 0 _053_
rlabel via2 78 36708 78 36708 0 clk
rlabel metal2 33216 22680 33216 22680 0 clknet_0_clk
rlabel metal3 17856 15540 17856 15540 0 clknet_2_0__leaf_clk
rlabel metal2 16224 23100 16224 23100 0 clknet_2_1__leaf_clk
rlabel metal3 39456 19236 39456 19236 0 clknet_2_2__leaf_clk
rlabel metal3 37872 23100 37872 23100 0 clknet_2_3__leaf_clk
rlabel metal2 28608 22974 28608 22974 0 mod1.bpsk_mod.i_out\[2\]
rlabel metal3 18048 15708 18048 15708 0 mod1.i_out_8psk\[0\]
rlabel metal2 28800 22302 28800 22302 0 mod1.i_out_8psk\[1\]
rlabel metal3 35952 22260 35952 22260 0 mod1.i_out_8psk\[2\]
rlabel metal2 32448 22176 32448 22176 0 mod1.i_out_qam16\[2\]
rlabel metal2 35808 22302 35808 22302 0 mod1.i_out_qam16\[3\]
rlabel metal2 39264 16254 39264 16254 0 mod1.i_out_qpsk\[1\]
rlabel metal3 37488 20076 37488 20076 0 mod1.i_out_qpsk\[2\]
rlabel metal2 33792 16926 33792 16926 0 mod1.psk8_mod.q_out\[1\]
rlabel metal3 26496 15540 26496 15540 0 mod1.psk8_mod.q_out\[2\]
rlabel metal2 26784 12390 26784 12390 0 mod1.q_out_qam16\[2\]
rlabel metal3 25680 11928 25680 11928 0 mod1.q_out_qam16\[3\]
rlabel metal2 29184 17724 29184 17724 0 mod1.q_out_qpsk\[2\]
rlabel metal2 14976 21168 14976 21168 0 mod1.qam16_mod.i_level\[2\]
rlabel metal2 22464 18606 22464 18606 0 mod1.qam16_mod.i_level\[3\]
rlabel metal2 17616 18648 17616 18648 0 mod1.qam16_mod.q_level\[2\]
rlabel metal2 21888 18060 21888 18060 0 mod1.qam16_mod.q_level\[3\]
rlabel metal3 15504 23772 15504 23772 0 net1
rlabel metal2 1056 29064 1056 29064 0 net10
rlabel metal2 35616 22344 35616 22344 0 net11
rlabel metal2 20448 26838 20448 26838 0 net12
rlabel metal2 37920 17430 37920 17430 0 net13
rlabel metal3 20832 23100 20832 23100 0 net14
rlabel metal2 39168 19152 39168 19152 0 net15
rlabel metal2 1152 30870 1152 30870 0 net16
rlabel metal3 14976 32844 14976 32844 0 net17
rlabel metal3 15264 33684 15264 33684 0 net18
rlabel metal3 15120 34356 15120 34356 0 net19
rlabel metal2 17760 19656 17760 19656 0 net2
rlabel metal2 23520 31668 23520 31668 0 net20
rlabel metal3 13968 9408 13968 9408 0 net21
rlabel metal2 36768 19950 36768 19950 0 net22
rlabel metal2 18048 13020 18048 13020 0 net23
rlabel metal2 864 12390 864 12390 0 net24
rlabel metal2 816 2688 816 2688 0 net25
rlabel metal2 1008 3360 1008 3360 0 net26
rlabel metal2 34464 13146 34464 13146 0 net27
rlabel metal3 34368 22008 34368 22008 0 net28
rlabel metal2 18912 15414 18912 15414 0 net29
rlabel metal2 18048 19026 18048 19026 0 net3
rlabel metal2 34272 12012 34272 12012 0 net30
rlabel metal2 1056 9954 1056 9954 0 net31
rlabel metal2 768 10458 768 10458 0 net32
rlabel metal3 366 12348 366 12348 0 net33
rlabel metal3 366 13188 366 13188 0 net34
rlabel metal3 366 14028 366 14028 0 net35
rlabel metal3 366 14868 366 14868 0 net36
rlabel metal2 30912 12432 30912 12432 0 net37
rlabel metal3 318 15708 318 15708 0 net38
rlabel metal3 366 16548 366 16548 0 net39
rlabel metal2 21264 20076 21264 20076 0 net4
rlabel metal3 366 17388 366 17388 0 net40
rlabel metal3 366 18228 366 18228 0 net41
rlabel metal3 366 19068 366 19068 0 net42
rlabel metal3 366 19908 366 19908 0 net43
rlabel metal3 366 20748 366 20748 0 net44
rlabel metal3 78 21588 78 21588 0 net45
rlabel metal3 37968 16212 37968 16212 0 net46
rlabel metal3 27936 18564 27936 18564 0 net47
rlabel metal2 37248 19530 37248 19530 0 net48
rlabel metal2 22560 17388 22560 17388 0 net5
rlabel metal2 960 26208 960 26208 0 net6
rlabel metal2 29184 20832 29184 20832 0 net7
rlabel metal2 960 28560 960 28560 0 net8
rlabel metal2 768 29106 768 29106 0 net9
rlabel metal3 174 37548 174 37548 0 rst_n
rlabel metal3 366 23268 366 23268 0 ui_in[1]
rlabel metal3 366 24108 366 24108 0 ui_in[2]
rlabel metal3 366 24948 366 24948 0 ui_in[3]
rlabel metal3 366 25788 366 25788 0 ui_in[4]
rlabel metal3 366 26628 366 26628 0 ui_in[5]
rlabel metal3 366 27468 366 27468 0 ui_in[6]
rlabel metal3 366 28308 366 28308 0 ui_in[7]
rlabel metal3 366 29148 366 29148 0 uio_in[0]
rlabel metal3 366 29988 366 29988 0 uio_in[1]
rlabel metal3 366 30828 366 30828 0 uio_in[2]
rlabel metal3 366 31668 366 31668 0 uio_in[3]
rlabel metal3 366 32508 366 32508 0 uio_in[4]
rlabel metal3 366 33348 366 33348 0 uio_in[5]
rlabel metal3 366 34188 366 34188 0 uio_in[6]
rlabel metal3 366 35028 366 35028 0 uio_in[7]
rlabel metal3 366 8988 366 8988 0 uio_out[0]
rlabel metal3 366 9828 366 9828 0 uio_out[1]
rlabel metal3 366 10668 366 10668 0 uio_out[2]
rlabel metal3 366 11508 366 11508 0 uio_out[3]
rlabel metal3 366 2268 366 2268 0 uo_out[0]
rlabel metal3 366 3108 366 3108 0 uo_out[1]
rlabel metal3 366 3948 366 3948 0 uo_out[2]
rlabel metal3 366 4788 366 4788 0 uo_out[3]
rlabel metal3 366 5628 366 5628 0 uo_out[4]
rlabel metal3 366 6468 366 6468 0 uo_out[5]
rlabel metal3 366 7308 366 7308 0 uo_out[6]
rlabel metal3 366 8148 366 8148 0 uo_out[7]
<< properties >>
string FIXED_BBOX 0 0 100000 40000
<< end >>
