module heichips25_template (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire \Demo1.epsk_de1.bit_out[0] ;
 wire \Demo1.epsk_de1.bit_out[1] ;
 wire \Demo1.epsk_de1.bit_out[2] ;
 wire \Demo1.qam16_bits[0] ;
 wire \Demo1.qam16_bits[1] ;
 wire \Demo1.qam16_bits[2] ;
 wire \Demo1.qam16_bits[3] ;
 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire net38;
 wire \mod1.bpsk_mod.i_out[2] ;
 wire \mod1.i_out_8psk[0] ;
 wire \mod1.i_out_8psk[1] ;
 wire \mod1.i_out_8psk[2] ;
 wire \mod1.i_out_qam16[2] ;
 wire \mod1.i_out_qam16[3] ;
 wire \mod1.i_out_qpsk[1] ;
 wire \mod1.i_out_qpsk[2] ;
 wire \mod1.psk8_mod.q_out[1] ;
 wire \mod1.psk8_mod.q_out[2] ;
 wire \mod1.q_out_qam16[2] ;
 wire \mod1.q_out_qam16[3] ;
 wire \mod1.q_out_qpsk[2] ;
 wire \mod1.qam16_mod.i_level[2] ;
 wire \mod1.qam16_mod.i_level[3] ;
 wire \mod1.qam16_mod.q_level[2] ;
 wire \mod1.qam16_mod.q_level[3] ;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire clknet_0_clk;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net33;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire net46;
 wire net47;
 wire net48;

 sg13g2_inv_1 _055_ (.Y(\mod1.qam16_mod.q_level[3] ),
    .A(net3));
 sg13g2_inv_1 _056_ (.Y(_032_),
    .A(net4));
 sg13g2_inv_4 _057_ (.A(net5),
    .Y(\mod1.qam16_mod.i_level[3] ));
 sg13g2_inv_1 _058_ (.Y(_033_),
    .A(net7));
 sg13g2_inv_1 _059_ (.Y(_034_),
    .A(net6));
 sg13g2_inv_1 _060_ (.Y(_035_),
    .A(net47));
 sg13g2_and2_1 _061_ (.A(net7),
    .B(net6),
    .X(_036_));
 sg13g2_or2_1 _062_ (.X(_037_),
    .B(net10),
    .A(net16));
 sg13g2_and2_1 _063_ (.A(net9),
    .B(net8),
    .X(_038_));
 sg13g2_o21ai_1 _064_ (.B1(net12),
    .Y(_011_),
    .A1(_037_),
    .A2(_038_));
 sg13g2_nand2_2 _065_ (.Y(_039_),
    .A(_032_),
    .B(\mod1.qam16_mod.i_level[3] ));
 sg13g2_nor2_2 _066_ (.A(net3),
    .B(net4),
    .Y(_040_));
 sg13g2_nand3b_1 _067_ (.B(\mod1.qam16_mod.i_level[3] ),
    .C(_040_),
    .Y(_000_),
    .A_N(net2));
 sg13g2_nor2b_2 _068_ (.A(net6),
    .B_N(net7),
    .Y(_041_));
 sg13g2_a22oi_1 _069_ (.Y(_042_),
    .B1(_041_),
    .B2(\Demo1.epsk_de1.bit_out[0] ),
    .A2(net11),
    .A1(\Demo1.qam16_bits[0] ));
 sg13g2_inv_4 _070_ (.A(_042_),
    .Y(net21));
 sg13g2_a22oi_1 _071_ (.Y(_043_),
    .B1(_041_),
    .B2(\Demo1.epsk_de1.bit_out[1] ),
    .A2(net11),
    .A1(\Demo1.qam16_bits[1] ));
 sg13g2_inv_4 _072_ (.A(_043_),
    .Y(net22));
 sg13g2_a22oi_1 _073_ (.Y(_044_),
    .B1(_041_),
    .B2(\Demo1.epsk_de1.bit_out[2] ),
    .A2(net12),
    .A1(\Demo1.qam16_bits[2] ));
 sg13g2_inv_2 _074_ (.Y(net23),
    .A(_044_));
 sg13g2_and2_1 _075_ (.A(\Demo1.qam16_bits[3] ),
    .B(net11),
    .X(net24));
 sg13g2_xor2_1 _076_ (.B(net5),
    .A(net4),
    .X(\mod1.qam16_mod.i_level[2] ));
 sg13g2_and2_1 _077_ (.A(\mod1.i_out_8psk[0] ),
    .B(_041_),
    .X(net29));
 sg13g2_nor2b_2 _078_ (.A(net7),
    .B_N(net6),
    .Y(_045_));
 sg13g2_a22oi_1 _079_ (.Y(_046_),
    .B1(_045_),
    .B2(\mod1.i_out_qpsk[1] ),
    .A2(net11),
    .A1(\Demo1.qam16_bits[3] ));
 sg13g2_o21ai_1 _080_ (.B1(_034_),
    .Y(_047_),
    .A1(_033_),
    .A2(\mod1.i_out_8psk[1] ));
 sg13g2_nor3_1 _081_ (.A(net7),
    .B(net6),
    .C(\Demo1.qam16_bits[3] ),
    .Y(_048_));
 sg13g2_a21oi_2 _082_ (.B1(_048_),
    .Y(net26),
    .A2(_047_),
    .A1(_046_));
 sg13g2_nand2_1 _083_ (.Y(_049_),
    .A(\mod1.i_out_8psk[2] ),
    .B(_041_));
 sg13g2_nand2_1 _084_ (.Y(_050_),
    .A(\mod1.i_out_qpsk[2] ),
    .B(_045_));
 sg13g2_nand3_1 _085_ (.B(_034_),
    .C(\mod1.bpsk_mod.i_out[2] ),
    .A(_033_),
    .Y(_051_));
 sg13g2_nand2_1 _086_ (.Y(_052_),
    .A(\mod1.i_out_qam16[2] ),
    .B(net11));
 sg13g2_nand4_1 _087_ (.B(_050_),
    .C(_051_),
    .A(_049_),
    .Y(net27),
    .D(_052_));
 sg13g2_nand2_1 _088_ (.Y(_053_),
    .A(\mod1.i_out_qam16[3] ),
    .B(net11));
 sg13g2_nand4_1 _089_ (.B(_050_),
    .C(_051_),
    .A(_049_),
    .Y(net28),
    .D(_053_));
 sg13g2_nand2_1 _090_ (.Y(_015_),
    .A(\mod1.psk8_mod.q_out[1] ),
    .B(_041_));
 sg13g2_nand2_2 _091_ (.Y(net30),
    .A(_046_),
    .B(_015_));
 sg13g2_a22oi_1 _092_ (.Y(_016_),
    .B1(_045_),
    .B2(\mod1.q_out_qpsk[2] ),
    .A2(_041_),
    .A1(\mod1.psk8_mod.q_out[2] ));
 sg13g2_nand2_1 _093_ (.Y(_017_),
    .A(\mod1.q_out_qam16[2] ),
    .B(net11));
 sg13g2_nand2_2 _094_ (.Y(net31),
    .A(_016_),
    .B(_017_));
 sg13g2_nand2_1 _095_ (.Y(_018_),
    .A(\mod1.q_out_qam16[3] ),
    .B(net11));
 sg13g2_nand2_2 _096_ (.Y(net32),
    .A(_016_),
    .B(_018_));
 sg13g2_nor2_1 _097_ (.A(\mod1.qam16_mod.q_level[3] ),
    .B(net2),
    .Y(_019_));
 sg13g2_nand2b_1 _098_ (.Y(_020_),
    .B(net3),
    .A_N(net2));
 sg13g2_xor2_1 _099_ (.B(net2),
    .A(net3),
    .X(\mod1.qam16_mod.q_level[2] ));
 sg13g2_xnor2_1 _100_ (.Y(_021_),
    .A(net4),
    .B(\mod1.qam16_mod.q_level[2] ));
 sg13g2_nor2_1 _101_ (.A(net5),
    .B(_021_),
    .Y(_006_));
 sg13g2_nand3_1 _102_ (.B(net4),
    .C(\mod1.qam16_mod.i_level[3] ),
    .A(net3),
    .Y(_022_));
 sg13g2_o21ai_1 _103_ (.B1(_022_),
    .Y(_007_),
    .A1(net2),
    .A2(_039_));
 sg13g2_o21ai_1 _104_ (.B1(_022_),
    .Y(_008_),
    .A1(_039_),
    .A2(_020_));
 sg13g2_nor3_1 _105_ (.A(net5),
    .B(_040_),
    .C(_019_),
    .Y(_009_));
 sg13g2_nor3_1 _106_ (.A(_032_),
    .B(net5),
    .C(_019_),
    .Y(_010_));
 sg13g2_and2_1 _107_ (.A(net20),
    .B(net12),
    .X(_023_));
 sg13g2_inv_1 _108_ (.Y(_005_),
    .A(_023_));
 sg13g2_or2_1 _109_ (.X(_024_),
    .B(net1),
    .A(net17));
 sg13g2_nand3_1 _110_ (.B(net18),
    .C(_024_),
    .A(net19),
    .Y(_025_));
 sg13g2_or2_1 _111_ (.X(_026_),
    .B(net18),
    .A(net19));
 sg13g2_a21o_1 _112_ (.A2(net1),
    .A1(net17),
    .B1(_026_),
    .X(_027_));
 sg13g2_nor2b_1 _113_ (.A(net20),
    .B_N(net12),
    .Y(_028_));
 sg13g2_a22oi_1 _114_ (.Y(_004_),
    .B1(_027_),
    .B2(_028_),
    .A2(_025_),
    .A1(_023_));
 sg13g2_nor4_1 _115_ (.A(net19),
    .B(net18),
    .C(net17),
    .D(net1),
    .Y(_029_));
 sg13g2_nor4_1 _116_ (.A(_033_),
    .B(net6),
    .C(net20),
    .D(_029_),
    .Y(_030_));
 sg13g2_and2_1 _117_ (.A(net20),
    .B(_041_),
    .X(_003_));
 sg13g2_nor3_1 _118_ (.A(net9),
    .B(net8),
    .C(_037_),
    .Y(_031_));
 sg13g2_a21o_1 _119_ (.A2(_031_),
    .A1(_003_),
    .B1(_030_),
    .X(_001_));
 sg13g2_and2_1 _120_ (.A(_030_),
    .B(_031_),
    .X(_002_));
 sg13g2_nand2b_1 _121_ (.Y(_012_),
    .B(_039_),
    .A_N(net46));
 sg13g2_mux2_1 _122_ (.A0(net2),
    .A1(net48),
    .S(_039_),
    .X(_013_));
 sg13g2_a22oi_1 _123_ (.Y(_014_),
    .B1(_040_),
    .B2(\mod1.qam16_mod.i_level[3] ),
    .A2(_039_),
    .A1(_035_));
 sg13g2_dfrbpq_1 _124_ (.RESET_B(net13),
    .D(\mod1.qam16_mod.q_level[2] ),
    .Q(\mod1.q_out_qam16[2] ),
    .CLK(clknet_2_0__leaf_clk));
 sg13g2_dfrbpq_1 _125_ (.RESET_B(net13),
    .D(\mod1.qam16_mod.q_level[3] ),
    .Q(\mod1.q_out_qam16[3] ),
    .CLK(clknet_2_0__leaf_clk));
 sg13g2_dfrbpq_1 _126_ (.RESET_B(net13),
    .D(_009_),
    .Q(\mod1.psk8_mod.q_out[1] ),
    .CLK(clknet_2_2__leaf_clk));
 sg13g2_dfrbpq_1 _127_ (.RESET_B(net13),
    .D(_010_),
    .Q(\mod1.psk8_mod.q_out[2] ),
    .CLK(clknet_2_0__leaf_clk));
 sg13g2_dfrbpq_1 _128_ (.RESET_B(net13),
    .D(_006_),
    .Q(\mod1.i_out_8psk[0] ),
    .CLK(clknet_2_0__leaf_clk));
 sg13g2_dfrbpq_1 _129_ (.RESET_B(net14),
    .D(_007_),
    .Q(\mod1.i_out_8psk[1] ),
    .CLK(clknet_2_3__leaf_clk));
 sg13g2_dfrbpq_1 _130_ (.RESET_B(net15),
    .D(_008_),
    .Q(\mod1.i_out_8psk[2] ),
    .CLK(clknet_2_3__leaf_clk));
 sg13g2_dfrbpq_1 _131_ (.RESET_B(net14),
    .D(\mod1.qam16_mod.i_level[2] ),
    .Q(\mod1.i_out_qam16[2] ),
    .CLK(clknet_2_1__leaf_clk));
 sg13g2_dfrbpq_1 _132_ (.RESET_B(net15),
    .D(\mod1.qam16_mod.i_level[3] ),
    .Q(\mod1.i_out_qam16[3] ),
    .CLK(clknet_2_3__leaf_clk));
 sg13g2_dfrbpq_1 _133_ (.RESET_B(net13),
    .D(_012_),
    .Q(\mod1.i_out_qpsk[1] ),
    .CLK(clknet_2_2__leaf_clk));
 sg13g2_dfrbpq_1 _134_ (.RESET_B(net15),
    .D(_013_),
    .Q(\mod1.i_out_qpsk[2] ),
    .CLK(clknet_2_2__leaf_clk));
 sg13g2_dfrbpq_1 _135_ (.RESET_B(net14),
    .D(_004_),
    .Q(\Demo1.qam16_bits[0] ),
    .CLK(clknet_2_1__leaf_clk));
 sg13g2_dfrbpq_1 _136_ (.RESET_B(net14),
    .D(_005_),
    .Q(\Demo1.qam16_bits[1] ),
    .CLK(clknet_2_3__leaf_clk));
 sg13g2_dfrbpq_1 _137_ (.RESET_B(net14),
    .D(_011_),
    .Q(\Demo1.qam16_bits[2] ),
    .CLK(clknet_2_1__leaf_clk));
 sg13g2_dfrbpq_1 _138_ (.RESET_B(net14),
    .D(_001_),
    .Q(\Demo1.epsk_de1.bit_out[0] ),
    .CLK(clknet_2_1__leaf_clk));
 sg13g2_dfrbpq_1 _139_ (.RESET_B(net15),
    .D(_002_),
    .Q(\Demo1.epsk_de1.bit_out[1] ),
    .CLK(clknet_2_3__leaf_clk));
 sg13g2_dfrbpq_1 _140_ (.RESET_B(net14),
    .D(_003_),
    .Q(\Demo1.epsk_de1.bit_out[2] ),
    .CLK(clknet_2_1__leaf_clk));
 sg13g2_dfrbpq_1 _141_ (.RESET_B(net13),
    .D(_014_),
    .Q(\mod1.q_out_qpsk[2] ),
    .CLK(clknet_2_2__leaf_clk));
 sg13g2_dfrbpq_2 _142_ (.RESET_B(net13),
    .D(net37),
    .Q(\Demo1.qam16_bits[3] ),
    .CLK(clknet_2_2__leaf_clk));
 sg13g2_dfrbpq_1 _143_ (.RESET_B(net14),
    .D(_000_),
    .Q(\mod1.bpsk_mod.i_out[2] ),
    .CLK(clknet_2_0__leaf_clk));
 sg13g2_tiehi heichips25_template_33 (.L_HI(net38));
 sg13g2_tiehi heichips25_template_34 (.L_HI(net39));
 sg13g2_tiehi heichips25_template_35 (.L_HI(net40));
 sg13g2_tiehi heichips25_template_36 (.L_HI(net41));
 sg13g2_tiehi heichips25_template_37 (.L_HI(net42));
 sg13g2_tiehi heichips25_template_38 (.L_HI(net43));
 sg13g2_tiehi heichips25_template_39 (.L_HI(net44));
 sg13g2_tiehi heichips25_template_40 (.L_HI(net45));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo heichips25_template_29 (.L_LO(net34));
 sg13g2_tielo heichips25_template_30 (.L_LO(net35));
 sg13g2_tielo heichips25_template_31 (.L_LO(net36));
 sg13g2_tiehi _142__32 (.L_HI(net37));
 sg13g2_buf_1 _157_ (.A(net29),
    .X(net25));
 sg13g2_buf_8 fanout11 (.A(_036_),
    .X(net11));
 sg13g2_buf_1 fanout12 (.A(_036_),
    .X(net12));
 sg13g2_buf_8 fanout13 (.A(net15),
    .X(net13));
 sg13g2_buf_8 fanout14 (.A(net15),
    .X(net14));
 sg13g2_buf_8 fanout15 (.A(rst_n),
    .X(net15));
 sg13g2_buf_2 input1 (.A(ui_in[1]),
    .X(net1));
 sg13g2_buf_2 input2 (.A(ui_in[2]),
    .X(net2));
 sg13g2_buf_2 input3 (.A(ui_in[3]),
    .X(net3));
 sg13g2_buf_2 input4 (.A(ui_in[4]),
    .X(net4));
 sg13g2_buf_2 input5 (.A(ui_in[5]),
    .X(net5));
 sg13g2_buf_2 input6 (.A(ui_in[6]),
    .X(net6));
 sg13g2_buf_2 input7 (.A(ui_in[7]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(uio_in[0]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(uio_in[1]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[2]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(uio_in[3]),
    .X(net16));
 sg13g2_buf_2 input12 (.A(uio_in[4]),
    .X(net17));
 sg13g2_buf_2 input13 (.A(uio_in[5]),
    .X(net18));
 sg13g2_buf_2 input14 (.A(uio_in[6]),
    .X(net19));
 sg13g2_buf_2 input15 (.A(uio_in[7]),
    .X(net20));
 sg13g2_buf_1 output16 (.A(net21),
    .X(uio_out[0]));
 sg13g2_buf_1 output17 (.A(net22),
    .X(uio_out[1]));
 sg13g2_buf_1 output18 (.A(net23),
    .X(uio_out[2]));
 sg13g2_buf_1 output19 (.A(net24),
    .X(uio_out[3]));
 sg13g2_buf_1 output20 (.A(net25),
    .X(uo_out[0]));
 sg13g2_buf_1 output21 (.A(net26),
    .X(uo_out[1]));
 sg13g2_buf_1 output22 (.A(net27),
    .X(uo_out[2]));
 sg13g2_buf_1 output23 (.A(net28),
    .X(uo_out[3]));
 sg13g2_buf_1 output24 (.A(net29),
    .X(uo_out[4]));
 sg13g2_buf_1 output25 (.A(net30),
    .X(uo_out[5]));
 sg13g2_buf_1 output26 (.A(net31),
    .X(uo_out[6]));
 sg13g2_buf_1 output27 (.A(net32),
    .X(uo_out[7]));
 sg13g2_tielo heichips25_template_28 (.L_LO(net33));
 sg13g2_buf_8 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sg13g2_buf_8 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sg13g2_buf_8 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sg13g2_buf_8 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sg13g2_buf_1 clkload0 (.A(clknet_2_0__leaf_clk));
 sg13g2_buf_1 clkload1 (.A(clknet_2_1__leaf_clk));
 sg13g2_buf_1 clkload2 (.A(clknet_2_3__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\mod1.i_out_qpsk[1] ),
    .X(net46));
 sg13g2_dlygate4sd3_1 hold2 (.A(\mod1.q_out_qpsk[2] ),
    .X(net47));
 sg13g2_dlygate4sd3_1 hold3 (.A(\mod1.i_out_qpsk[2] ),
    .X(net48));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_decap_8 FILLER_0_427 ();
 sg13g2_decap_8 FILLER_0_434 ();
 sg13g2_decap_8 FILLER_0_441 ();
 sg13g2_decap_8 FILLER_0_448 ();
 sg13g2_decap_8 FILLER_0_455 ();
 sg13g2_decap_8 FILLER_0_462 ();
 sg13g2_decap_8 FILLER_0_469 ();
 sg13g2_decap_8 FILLER_0_476 ();
 sg13g2_decap_8 FILLER_0_483 ();
 sg13g2_decap_8 FILLER_0_490 ();
 sg13g2_decap_8 FILLER_0_497 ();
 sg13g2_decap_8 FILLER_0_504 ();
 sg13g2_decap_8 FILLER_0_511 ();
 sg13g2_decap_8 FILLER_0_518 ();
 sg13g2_decap_8 FILLER_0_525 ();
 sg13g2_decap_8 FILLER_0_532 ();
 sg13g2_decap_8 FILLER_0_539 ();
 sg13g2_decap_8 FILLER_0_546 ();
 sg13g2_decap_8 FILLER_0_553 ();
 sg13g2_decap_8 FILLER_0_560 ();
 sg13g2_decap_8 FILLER_0_567 ();
 sg13g2_decap_8 FILLER_0_574 ();
 sg13g2_decap_8 FILLER_0_581 ();
 sg13g2_decap_8 FILLER_0_588 ();
 sg13g2_decap_8 FILLER_0_595 ();
 sg13g2_decap_8 FILLER_0_602 ();
 sg13g2_decap_8 FILLER_0_609 ();
 sg13g2_decap_8 FILLER_0_616 ();
 sg13g2_decap_8 FILLER_0_623 ();
 sg13g2_decap_8 FILLER_0_630 ();
 sg13g2_decap_8 FILLER_0_637 ();
 sg13g2_decap_8 FILLER_0_644 ();
 sg13g2_decap_8 FILLER_0_651 ();
 sg13g2_decap_8 FILLER_0_658 ();
 sg13g2_decap_8 FILLER_0_665 ();
 sg13g2_decap_8 FILLER_0_672 ();
 sg13g2_decap_8 FILLER_0_679 ();
 sg13g2_decap_8 FILLER_0_686 ();
 sg13g2_decap_8 FILLER_0_693 ();
 sg13g2_decap_8 FILLER_0_700 ();
 sg13g2_decap_8 FILLER_0_707 ();
 sg13g2_decap_8 FILLER_0_714 ();
 sg13g2_decap_8 FILLER_0_721 ();
 sg13g2_decap_8 FILLER_0_728 ();
 sg13g2_decap_8 FILLER_0_735 ();
 sg13g2_decap_8 FILLER_0_742 ();
 sg13g2_decap_8 FILLER_0_749 ();
 sg13g2_decap_8 FILLER_0_756 ();
 sg13g2_decap_8 FILLER_0_763 ();
 sg13g2_decap_8 FILLER_0_770 ();
 sg13g2_decap_8 FILLER_0_777 ();
 sg13g2_decap_8 FILLER_0_784 ();
 sg13g2_decap_8 FILLER_0_791 ();
 sg13g2_decap_8 FILLER_0_798 ();
 sg13g2_decap_8 FILLER_0_805 ();
 sg13g2_decap_8 FILLER_0_812 ();
 sg13g2_decap_8 FILLER_0_819 ();
 sg13g2_decap_8 FILLER_0_826 ();
 sg13g2_decap_8 FILLER_0_833 ();
 sg13g2_decap_8 FILLER_0_840 ();
 sg13g2_decap_8 FILLER_0_847 ();
 sg13g2_decap_8 FILLER_0_854 ();
 sg13g2_decap_8 FILLER_0_861 ();
 sg13g2_decap_8 FILLER_0_868 ();
 sg13g2_decap_8 FILLER_0_875 ();
 sg13g2_decap_8 FILLER_0_882 ();
 sg13g2_decap_8 FILLER_0_889 ();
 sg13g2_decap_8 FILLER_0_896 ();
 sg13g2_decap_8 FILLER_0_903 ();
 sg13g2_decap_8 FILLER_0_910 ();
 sg13g2_decap_8 FILLER_0_917 ();
 sg13g2_decap_8 FILLER_0_924 ();
 sg13g2_decap_8 FILLER_0_931 ();
 sg13g2_decap_8 FILLER_0_938 ();
 sg13g2_decap_8 FILLER_0_945 ();
 sg13g2_decap_8 FILLER_0_952 ();
 sg13g2_decap_8 FILLER_0_959 ();
 sg13g2_decap_8 FILLER_0_966 ();
 sg13g2_decap_8 FILLER_0_973 ();
 sg13g2_decap_8 FILLER_0_980 ();
 sg13g2_decap_8 FILLER_0_987 ();
 sg13g2_decap_8 FILLER_0_994 ();
 sg13g2_decap_8 FILLER_0_1001 ();
 sg13g2_decap_8 FILLER_0_1008 ();
 sg13g2_decap_8 FILLER_0_1015 ();
 sg13g2_decap_8 FILLER_0_1022 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_decap_8 FILLER_1_427 ();
 sg13g2_decap_8 FILLER_1_434 ();
 sg13g2_decap_8 FILLER_1_441 ();
 sg13g2_decap_8 FILLER_1_448 ();
 sg13g2_decap_8 FILLER_1_455 ();
 sg13g2_decap_8 FILLER_1_462 ();
 sg13g2_decap_8 FILLER_1_469 ();
 sg13g2_decap_8 FILLER_1_476 ();
 sg13g2_decap_8 FILLER_1_483 ();
 sg13g2_decap_8 FILLER_1_490 ();
 sg13g2_decap_8 FILLER_1_497 ();
 sg13g2_decap_8 FILLER_1_504 ();
 sg13g2_decap_8 FILLER_1_511 ();
 sg13g2_decap_8 FILLER_1_518 ();
 sg13g2_decap_8 FILLER_1_525 ();
 sg13g2_decap_8 FILLER_1_532 ();
 sg13g2_decap_8 FILLER_1_539 ();
 sg13g2_decap_8 FILLER_1_546 ();
 sg13g2_decap_8 FILLER_1_553 ();
 sg13g2_decap_8 FILLER_1_560 ();
 sg13g2_decap_8 FILLER_1_567 ();
 sg13g2_decap_8 FILLER_1_574 ();
 sg13g2_decap_8 FILLER_1_581 ();
 sg13g2_decap_8 FILLER_1_588 ();
 sg13g2_decap_8 FILLER_1_595 ();
 sg13g2_decap_8 FILLER_1_602 ();
 sg13g2_decap_8 FILLER_1_609 ();
 sg13g2_decap_8 FILLER_1_616 ();
 sg13g2_decap_8 FILLER_1_623 ();
 sg13g2_decap_8 FILLER_1_630 ();
 sg13g2_decap_8 FILLER_1_637 ();
 sg13g2_decap_8 FILLER_1_644 ();
 sg13g2_decap_8 FILLER_1_651 ();
 sg13g2_decap_8 FILLER_1_658 ();
 sg13g2_decap_8 FILLER_1_665 ();
 sg13g2_decap_8 FILLER_1_672 ();
 sg13g2_decap_8 FILLER_1_679 ();
 sg13g2_decap_8 FILLER_1_686 ();
 sg13g2_decap_8 FILLER_1_693 ();
 sg13g2_decap_8 FILLER_1_700 ();
 sg13g2_decap_8 FILLER_1_707 ();
 sg13g2_decap_8 FILLER_1_714 ();
 sg13g2_decap_8 FILLER_1_721 ();
 sg13g2_decap_8 FILLER_1_728 ();
 sg13g2_decap_8 FILLER_1_735 ();
 sg13g2_decap_8 FILLER_1_742 ();
 sg13g2_decap_8 FILLER_1_749 ();
 sg13g2_decap_8 FILLER_1_756 ();
 sg13g2_decap_8 FILLER_1_763 ();
 sg13g2_decap_8 FILLER_1_770 ();
 sg13g2_decap_8 FILLER_1_777 ();
 sg13g2_decap_8 FILLER_1_784 ();
 sg13g2_decap_8 FILLER_1_791 ();
 sg13g2_decap_8 FILLER_1_798 ();
 sg13g2_decap_8 FILLER_1_805 ();
 sg13g2_decap_8 FILLER_1_812 ();
 sg13g2_decap_8 FILLER_1_819 ();
 sg13g2_decap_8 FILLER_1_826 ();
 sg13g2_decap_8 FILLER_1_833 ();
 sg13g2_decap_8 FILLER_1_840 ();
 sg13g2_decap_8 FILLER_1_847 ();
 sg13g2_decap_8 FILLER_1_854 ();
 sg13g2_decap_8 FILLER_1_861 ();
 sg13g2_decap_8 FILLER_1_868 ();
 sg13g2_decap_8 FILLER_1_875 ();
 sg13g2_decap_8 FILLER_1_882 ();
 sg13g2_decap_8 FILLER_1_889 ();
 sg13g2_decap_8 FILLER_1_896 ();
 sg13g2_decap_8 FILLER_1_903 ();
 sg13g2_decap_8 FILLER_1_910 ();
 sg13g2_decap_8 FILLER_1_917 ();
 sg13g2_decap_8 FILLER_1_924 ();
 sg13g2_decap_8 FILLER_1_931 ();
 sg13g2_decap_8 FILLER_1_938 ();
 sg13g2_decap_8 FILLER_1_945 ();
 sg13g2_decap_8 FILLER_1_952 ();
 sg13g2_decap_8 FILLER_1_959 ();
 sg13g2_decap_8 FILLER_1_966 ();
 sg13g2_decap_8 FILLER_1_973 ();
 sg13g2_decap_8 FILLER_1_980 ();
 sg13g2_decap_8 FILLER_1_987 ();
 sg13g2_decap_8 FILLER_1_994 ();
 sg13g2_decap_8 FILLER_1_1001 ();
 sg13g2_decap_8 FILLER_1_1008 ();
 sg13g2_decap_8 FILLER_1_1015 ();
 sg13g2_decap_8 FILLER_1_1022 ();
 sg13g2_decap_8 FILLER_2_4 ();
 sg13g2_decap_8 FILLER_2_11 ();
 sg13g2_decap_8 FILLER_2_18 ();
 sg13g2_decap_8 FILLER_2_25 ();
 sg13g2_decap_8 FILLER_2_32 ();
 sg13g2_decap_8 FILLER_2_39 ();
 sg13g2_decap_8 FILLER_2_46 ();
 sg13g2_decap_8 FILLER_2_53 ();
 sg13g2_decap_8 FILLER_2_60 ();
 sg13g2_decap_8 FILLER_2_67 ();
 sg13g2_decap_8 FILLER_2_74 ();
 sg13g2_decap_8 FILLER_2_81 ();
 sg13g2_decap_8 FILLER_2_88 ();
 sg13g2_decap_8 FILLER_2_95 ();
 sg13g2_decap_8 FILLER_2_102 ();
 sg13g2_decap_8 FILLER_2_109 ();
 sg13g2_decap_8 FILLER_2_116 ();
 sg13g2_decap_8 FILLER_2_123 ();
 sg13g2_decap_8 FILLER_2_130 ();
 sg13g2_decap_8 FILLER_2_137 ();
 sg13g2_decap_8 FILLER_2_144 ();
 sg13g2_decap_8 FILLER_2_151 ();
 sg13g2_decap_8 FILLER_2_158 ();
 sg13g2_decap_8 FILLER_2_165 ();
 sg13g2_decap_8 FILLER_2_172 ();
 sg13g2_decap_8 FILLER_2_179 ();
 sg13g2_decap_8 FILLER_2_186 ();
 sg13g2_decap_8 FILLER_2_193 ();
 sg13g2_decap_8 FILLER_2_200 ();
 sg13g2_decap_8 FILLER_2_207 ();
 sg13g2_decap_8 FILLER_2_214 ();
 sg13g2_decap_8 FILLER_2_221 ();
 sg13g2_decap_8 FILLER_2_228 ();
 sg13g2_decap_8 FILLER_2_235 ();
 sg13g2_decap_8 FILLER_2_242 ();
 sg13g2_decap_8 FILLER_2_249 ();
 sg13g2_decap_8 FILLER_2_256 ();
 sg13g2_decap_8 FILLER_2_263 ();
 sg13g2_decap_8 FILLER_2_270 ();
 sg13g2_decap_8 FILLER_2_277 ();
 sg13g2_decap_8 FILLER_2_284 ();
 sg13g2_decap_8 FILLER_2_291 ();
 sg13g2_decap_8 FILLER_2_298 ();
 sg13g2_decap_8 FILLER_2_305 ();
 sg13g2_decap_8 FILLER_2_312 ();
 sg13g2_decap_8 FILLER_2_319 ();
 sg13g2_decap_8 FILLER_2_326 ();
 sg13g2_decap_8 FILLER_2_333 ();
 sg13g2_decap_8 FILLER_2_340 ();
 sg13g2_decap_8 FILLER_2_347 ();
 sg13g2_decap_8 FILLER_2_354 ();
 sg13g2_decap_8 FILLER_2_361 ();
 sg13g2_decap_8 FILLER_2_368 ();
 sg13g2_decap_8 FILLER_2_375 ();
 sg13g2_decap_8 FILLER_2_382 ();
 sg13g2_decap_8 FILLER_2_389 ();
 sg13g2_decap_8 FILLER_2_396 ();
 sg13g2_decap_8 FILLER_2_403 ();
 sg13g2_decap_8 FILLER_2_410 ();
 sg13g2_decap_8 FILLER_2_417 ();
 sg13g2_decap_8 FILLER_2_424 ();
 sg13g2_decap_8 FILLER_2_431 ();
 sg13g2_decap_8 FILLER_2_438 ();
 sg13g2_decap_8 FILLER_2_445 ();
 sg13g2_decap_8 FILLER_2_452 ();
 sg13g2_decap_8 FILLER_2_459 ();
 sg13g2_decap_8 FILLER_2_466 ();
 sg13g2_decap_8 FILLER_2_473 ();
 sg13g2_decap_8 FILLER_2_480 ();
 sg13g2_decap_8 FILLER_2_487 ();
 sg13g2_decap_8 FILLER_2_494 ();
 sg13g2_decap_8 FILLER_2_501 ();
 sg13g2_decap_8 FILLER_2_508 ();
 sg13g2_decap_8 FILLER_2_515 ();
 sg13g2_decap_8 FILLER_2_522 ();
 sg13g2_decap_8 FILLER_2_529 ();
 sg13g2_decap_8 FILLER_2_536 ();
 sg13g2_decap_8 FILLER_2_543 ();
 sg13g2_decap_8 FILLER_2_550 ();
 sg13g2_decap_8 FILLER_2_557 ();
 sg13g2_decap_8 FILLER_2_564 ();
 sg13g2_decap_8 FILLER_2_571 ();
 sg13g2_decap_8 FILLER_2_578 ();
 sg13g2_decap_8 FILLER_2_585 ();
 sg13g2_decap_8 FILLER_2_592 ();
 sg13g2_decap_8 FILLER_2_599 ();
 sg13g2_decap_8 FILLER_2_606 ();
 sg13g2_decap_8 FILLER_2_613 ();
 sg13g2_decap_8 FILLER_2_620 ();
 sg13g2_decap_8 FILLER_2_627 ();
 sg13g2_decap_8 FILLER_2_634 ();
 sg13g2_decap_8 FILLER_2_641 ();
 sg13g2_decap_8 FILLER_2_648 ();
 sg13g2_decap_8 FILLER_2_655 ();
 sg13g2_decap_8 FILLER_2_662 ();
 sg13g2_decap_8 FILLER_2_669 ();
 sg13g2_decap_8 FILLER_2_676 ();
 sg13g2_decap_8 FILLER_2_683 ();
 sg13g2_decap_8 FILLER_2_690 ();
 sg13g2_decap_8 FILLER_2_697 ();
 sg13g2_decap_8 FILLER_2_704 ();
 sg13g2_decap_8 FILLER_2_711 ();
 sg13g2_decap_8 FILLER_2_718 ();
 sg13g2_decap_8 FILLER_2_725 ();
 sg13g2_decap_8 FILLER_2_732 ();
 sg13g2_decap_8 FILLER_2_739 ();
 sg13g2_decap_8 FILLER_2_746 ();
 sg13g2_decap_8 FILLER_2_753 ();
 sg13g2_decap_8 FILLER_2_760 ();
 sg13g2_decap_8 FILLER_2_767 ();
 sg13g2_decap_8 FILLER_2_774 ();
 sg13g2_decap_8 FILLER_2_781 ();
 sg13g2_decap_8 FILLER_2_788 ();
 sg13g2_decap_8 FILLER_2_795 ();
 sg13g2_decap_8 FILLER_2_802 ();
 sg13g2_decap_8 FILLER_2_809 ();
 sg13g2_decap_8 FILLER_2_816 ();
 sg13g2_decap_8 FILLER_2_823 ();
 sg13g2_decap_8 FILLER_2_830 ();
 sg13g2_decap_8 FILLER_2_837 ();
 sg13g2_decap_8 FILLER_2_844 ();
 sg13g2_decap_8 FILLER_2_851 ();
 sg13g2_decap_8 FILLER_2_858 ();
 sg13g2_decap_8 FILLER_2_865 ();
 sg13g2_decap_8 FILLER_2_872 ();
 sg13g2_decap_8 FILLER_2_879 ();
 sg13g2_decap_8 FILLER_2_886 ();
 sg13g2_decap_8 FILLER_2_893 ();
 sg13g2_decap_8 FILLER_2_900 ();
 sg13g2_decap_8 FILLER_2_907 ();
 sg13g2_decap_8 FILLER_2_914 ();
 sg13g2_decap_8 FILLER_2_921 ();
 sg13g2_decap_8 FILLER_2_928 ();
 sg13g2_decap_8 FILLER_2_935 ();
 sg13g2_decap_8 FILLER_2_942 ();
 sg13g2_decap_8 FILLER_2_949 ();
 sg13g2_decap_8 FILLER_2_956 ();
 sg13g2_decap_8 FILLER_2_963 ();
 sg13g2_decap_8 FILLER_2_970 ();
 sg13g2_decap_8 FILLER_2_977 ();
 sg13g2_decap_8 FILLER_2_984 ();
 sg13g2_decap_8 FILLER_2_991 ();
 sg13g2_decap_8 FILLER_2_998 ();
 sg13g2_decap_8 FILLER_2_1005 ();
 sg13g2_decap_8 FILLER_2_1012 ();
 sg13g2_decap_8 FILLER_2_1019 ();
 sg13g2_fill_2 FILLER_2_1026 ();
 sg13g2_fill_1 FILLER_2_1028 ();
 sg13g2_decap_8 FILLER_3_4 ();
 sg13g2_decap_8 FILLER_3_11 ();
 sg13g2_decap_8 FILLER_3_18 ();
 sg13g2_decap_8 FILLER_3_25 ();
 sg13g2_decap_8 FILLER_3_32 ();
 sg13g2_decap_8 FILLER_3_39 ();
 sg13g2_decap_8 FILLER_3_46 ();
 sg13g2_decap_8 FILLER_3_53 ();
 sg13g2_decap_8 FILLER_3_60 ();
 sg13g2_decap_8 FILLER_3_67 ();
 sg13g2_decap_8 FILLER_3_74 ();
 sg13g2_decap_8 FILLER_3_81 ();
 sg13g2_decap_8 FILLER_3_88 ();
 sg13g2_decap_8 FILLER_3_95 ();
 sg13g2_decap_8 FILLER_3_102 ();
 sg13g2_decap_8 FILLER_3_109 ();
 sg13g2_decap_8 FILLER_3_116 ();
 sg13g2_decap_8 FILLER_3_123 ();
 sg13g2_decap_8 FILLER_3_130 ();
 sg13g2_decap_8 FILLER_3_137 ();
 sg13g2_decap_8 FILLER_3_144 ();
 sg13g2_decap_8 FILLER_3_151 ();
 sg13g2_decap_8 FILLER_3_158 ();
 sg13g2_decap_8 FILLER_3_165 ();
 sg13g2_decap_8 FILLER_3_172 ();
 sg13g2_decap_8 FILLER_3_179 ();
 sg13g2_decap_8 FILLER_3_186 ();
 sg13g2_decap_8 FILLER_3_193 ();
 sg13g2_decap_8 FILLER_3_200 ();
 sg13g2_decap_8 FILLER_3_207 ();
 sg13g2_decap_8 FILLER_3_214 ();
 sg13g2_decap_8 FILLER_3_221 ();
 sg13g2_decap_8 FILLER_3_228 ();
 sg13g2_decap_8 FILLER_3_235 ();
 sg13g2_decap_8 FILLER_3_242 ();
 sg13g2_decap_8 FILLER_3_249 ();
 sg13g2_decap_8 FILLER_3_256 ();
 sg13g2_decap_8 FILLER_3_263 ();
 sg13g2_decap_8 FILLER_3_270 ();
 sg13g2_decap_8 FILLER_3_277 ();
 sg13g2_decap_8 FILLER_3_284 ();
 sg13g2_decap_8 FILLER_3_291 ();
 sg13g2_decap_8 FILLER_3_298 ();
 sg13g2_decap_8 FILLER_3_305 ();
 sg13g2_decap_8 FILLER_3_312 ();
 sg13g2_decap_8 FILLER_3_319 ();
 sg13g2_decap_8 FILLER_3_326 ();
 sg13g2_decap_8 FILLER_3_333 ();
 sg13g2_decap_8 FILLER_3_340 ();
 sg13g2_decap_8 FILLER_3_347 ();
 sg13g2_decap_8 FILLER_3_354 ();
 sg13g2_decap_8 FILLER_3_361 ();
 sg13g2_decap_8 FILLER_3_368 ();
 sg13g2_decap_8 FILLER_3_375 ();
 sg13g2_decap_8 FILLER_3_382 ();
 sg13g2_decap_8 FILLER_3_389 ();
 sg13g2_decap_8 FILLER_3_396 ();
 sg13g2_decap_8 FILLER_3_403 ();
 sg13g2_decap_8 FILLER_3_410 ();
 sg13g2_decap_8 FILLER_3_417 ();
 sg13g2_decap_8 FILLER_3_424 ();
 sg13g2_decap_8 FILLER_3_431 ();
 sg13g2_decap_8 FILLER_3_438 ();
 sg13g2_decap_8 FILLER_3_445 ();
 sg13g2_decap_8 FILLER_3_452 ();
 sg13g2_decap_8 FILLER_3_459 ();
 sg13g2_decap_8 FILLER_3_466 ();
 sg13g2_decap_8 FILLER_3_473 ();
 sg13g2_decap_8 FILLER_3_480 ();
 sg13g2_decap_8 FILLER_3_487 ();
 sg13g2_decap_8 FILLER_3_494 ();
 sg13g2_decap_8 FILLER_3_501 ();
 sg13g2_decap_8 FILLER_3_508 ();
 sg13g2_decap_8 FILLER_3_515 ();
 sg13g2_decap_8 FILLER_3_522 ();
 sg13g2_decap_8 FILLER_3_529 ();
 sg13g2_decap_8 FILLER_3_536 ();
 sg13g2_decap_8 FILLER_3_543 ();
 sg13g2_decap_8 FILLER_3_550 ();
 sg13g2_decap_8 FILLER_3_557 ();
 sg13g2_decap_8 FILLER_3_564 ();
 sg13g2_decap_8 FILLER_3_571 ();
 sg13g2_decap_8 FILLER_3_578 ();
 sg13g2_decap_8 FILLER_3_585 ();
 sg13g2_decap_8 FILLER_3_592 ();
 sg13g2_decap_8 FILLER_3_599 ();
 sg13g2_decap_8 FILLER_3_606 ();
 sg13g2_decap_8 FILLER_3_613 ();
 sg13g2_decap_8 FILLER_3_620 ();
 sg13g2_decap_8 FILLER_3_627 ();
 sg13g2_decap_8 FILLER_3_634 ();
 sg13g2_decap_8 FILLER_3_641 ();
 sg13g2_decap_8 FILLER_3_648 ();
 sg13g2_decap_8 FILLER_3_655 ();
 sg13g2_decap_8 FILLER_3_662 ();
 sg13g2_decap_8 FILLER_3_669 ();
 sg13g2_decap_8 FILLER_3_676 ();
 sg13g2_decap_8 FILLER_3_683 ();
 sg13g2_decap_8 FILLER_3_690 ();
 sg13g2_decap_8 FILLER_3_697 ();
 sg13g2_decap_8 FILLER_3_704 ();
 sg13g2_decap_8 FILLER_3_711 ();
 sg13g2_decap_8 FILLER_3_718 ();
 sg13g2_decap_8 FILLER_3_725 ();
 sg13g2_decap_8 FILLER_3_732 ();
 sg13g2_decap_8 FILLER_3_739 ();
 sg13g2_decap_8 FILLER_3_746 ();
 sg13g2_decap_8 FILLER_3_753 ();
 sg13g2_decap_8 FILLER_3_760 ();
 sg13g2_decap_8 FILLER_3_767 ();
 sg13g2_decap_8 FILLER_3_774 ();
 sg13g2_decap_8 FILLER_3_781 ();
 sg13g2_decap_8 FILLER_3_788 ();
 sg13g2_decap_8 FILLER_3_795 ();
 sg13g2_decap_8 FILLER_3_802 ();
 sg13g2_decap_8 FILLER_3_809 ();
 sg13g2_decap_8 FILLER_3_816 ();
 sg13g2_decap_8 FILLER_3_823 ();
 sg13g2_decap_8 FILLER_3_830 ();
 sg13g2_decap_8 FILLER_3_837 ();
 sg13g2_decap_8 FILLER_3_844 ();
 sg13g2_decap_8 FILLER_3_851 ();
 sg13g2_decap_8 FILLER_3_858 ();
 sg13g2_decap_8 FILLER_3_865 ();
 sg13g2_decap_8 FILLER_3_872 ();
 sg13g2_decap_8 FILLER_3_879 ();
 sg13g2_decap_8 FILLER_3_886 ();
 sg13g2_decap_8 FILLER_3_893 ();
 sg13g2_decap_8 FILLER_3_900 ();
 sg13g2_decap_8 FILLER_3_907 ();
 sg13g2_decap_8 FILLER_3_914 ();
 sg13g2_decap_8 FILLER_3_921 ();
 sg13g2_decap_8 FILLER_3_928 ();
 sg13g2_decap_8 FILLER_3_935 ();
 sg13g2_decap_8 FILLER_3_942 ();
 sg13g2_decap_8 FILLER_3_949 ();
 sg13g2_decap_8 FILLER_3_956 ();
 sg13g2_decap_8 FILLER_3_963 ();
 sg13g2_decap_8 FILLER_3_970 ();
 sg13g2_decap_8 FILLER_3_977 ();
 sg13g2_decap_8 FILLER_3_984 ();
 sg13g2_decap_8 FILLER_3_991 ();
 sg13g2_decap_8 FILLER_3_998 ();
 sg13g2_decap_8 FILLER_3_1005 ();
 sg13g2_decap_8 FILLER_3_1012 ();
 sg13g2_decap_8 FILLER_3_1019 ();
 sg13g2_fill_2 FILLER_3_1026 ();
 sg13g2_fill_1 FILLER_3_1028 ();
 sg13g2_decap_8 FILLER_4_4 ();
 sg13g2_decap_8 FILLER_4_11 ();
 sg13g2_decap_8 FILLER_4_18 ();
 sg13g2_decap_8 FILLER_4_25 ();
 sg13g2_decap_8 FILLER_4_32 ();
 sg13g2_decap_8 FILLER_4_39 ();
 sg13g2_decap_8 FILLER_4_46 ();
 sg13g2_decap_8 FILLER_4_53 ();
 sg13g2_decap_8 FILLER_4_60 ();
 sg13g2_decap_8 FILLER_4_67 ();
 sg13g2_decap_8 FILLER_4_74 ();
 sg13g2_decap_8 FILLER_4_81 ();
 sg13g2_decap_8 FILLER_4_88 ();
 sg13g2_decap_8 FILLER_4_95 ();
 sg13g2_decap_8 FILLER_4_102 ();
 sg13g2_decap_8 FILLER_4_109 ();
 sg13g2_decap_8 FILLER_4_116 ();
 sg13g2_decap_8 FILLER_4_123 ();
 sg13g2_decap_8 FILLER_4_130 ();
 sg13g2_decap_8 FILLER_4_137 ();
 sg13g2_decap_8 FILLER_4_144 ();
 sg13g2_decap_8 FILLER_4_151 ();
 sg13g2_decap_8 FILLER_4_158 ();
 sg13g2_decap_8 FILLER_4_165 ();
 sg13g2_decap_8 FILLER_4_172 ();
 sg13g2_decap_8 FILLER_4_179 ();
 sg13g2_decap_8 FILLER_4_186 ();
 sg13g2_decap_8 FILLER_4_193 ();
 sg13g2_decap_8 FILLER_4_200 ();
 sg13g2_decap_8 FILLER_4_207 ();
 sg13g2_decap_8 FILLER_4_214 ();
 sg13g2_decap_8 FILLER_4_221 ();
 sg13g2_decap_8 FILLER_4_228 ();
 sg13g2_decap_8 FILLER_4_235 ();
 sg13g2_decap_8 FILLER_4_242 ();
 sg13g2_decap_8 FILLER_4_249 ();
 sg13g2_decap_8 FILLER_4_256 ();
 sg13g2_decap_8 FILLER_4_263 ();
 sg13g2_decap_8 FILLER_4_270 ();
 sg13g2_decap_8 FILLER_4_277 ();
 sg13g2_decap_8 FILLER_4_284 ();
 sg13g2_decap_8 FILLER_4_291 ();
 sg13g2_decap_8 FILLER_4_298 ();
 sg13g2_decap_8 FILLER_4_305 ();
 sg13g2_decap_8 FILLER_4_312 ();
 sg13g2_decap_8 FILLER_4_319 ();
 sg13g2_decap_8 FILLER_4_326 ();
 sg13g2_decap_8 FILLER_4_333 ();
 sg13g2_decap_8 FILLER_4_340 ();
 sg13g2_decap_8 FILLER_4_347 ();
 sg13g2_decap_8 FILLER_4_354 ();
 sg13g2_decap_8 FILLER_4_361 ();
 sg13g2_decap_8 FILLER_4_368 ();
 sg13g2_decap_8 FILLER_4_375 ();
 sg13g2_decap_8 FILLER_4_382 ();
 sg13g2_decap_8 FILLER_4_389 ();
 sg13g2_decap_8 FILLER_4_396 ();
 sg13g2_decap_8 FILLER_4_403 ();
 sg13g2_decap_8 FILLER_4_410 ();
 sg13g2_decap_8 FILLER_4_417 ();
 sg13g2_decap_8 FILLER_4_424 ();
 sg13g2_decap_8 FILLER_4_431 ();
 sg13g2_decap_8 FILLER_4_438 ();
 sg13g2_decap_8 FILLER_4_445 ();
 sg13g2_decap_8 FILLER_4_452 ();
 sg13g2_decap_8 FILLER_4_459 ();
 sg13g2_decap_8 FILLER_4_466 ();
 sg13g2_decap_8 FILLER_4_473 ();
 sg13g2_decap_8 FILLER_4_480 ();
 sg13g2_decap_8 FILLER_4_487 ();
 sg13g2_decap_8 FILLER_4_494 ();
 sg13g2_decap_8 FILLER_4_501 ();
 sg13g2_decap_8 FILLER_4_508 ();
 sg13g2_decap_8 FILLER_4_515 ();
 sg13g2_decap_8 FILLER_4_522 ();
 sg13g2_decap_8 FILLER_4_529 ();
 sg13g2_decap_8 FILLER_4_536 ();
 sg13g2_decap_8 FILLER_4_543 ();
 sg13g2_decap_8 FILLER_4_550 ();
 sg13g2_decap_8 FILLER_4_557 ();
 sg13g2_decap_8 FILLER_4_564 ();
 sg13g2_decap_8 FILLER_4_571 ();
 sg13g2_decap_8 FILLER_4_578 ();
 sg13g2_decap_8 FILLER_4_585 ();
 sg13g2_decap_8 FILLER_4_592 ();
 sg13g2_decap_8 FILLER_4_599 ();
 sg13g2_decap_8 FILLER_4_606 ();
 sg13g2_decap_8 FILLER_4_613 ();
 sg13g2_decap_8 FILLER_4_620 ();
 sg13g2_decap_8 FILLER_4_627 ();
 sg13g2_decap_8 FILLER_4_634 ();
 sg13g2_decap_8 FILLER_4_641 ();
 sg13g2_decap_8 FILLER_4_648 ();
 sg13g2_decap_8 FILLER_4_655 ();
 sg13g2_decap_8 FILLER_4_662 ();
 sg13g2_decap_8 FILLER_4_669 ();
 sg13g2_decap_8 FILLER_4_676 ();
 sg13g2_decap_8 FILLER_4_683 ();
 sg13g2_decap_8 FILLER_4_690 ();
 sg13g2_decap_8 FILLER_4_697 ();
 sg13g2_decap_8 FILLER_4_704 ();
 sg13g2_decap_8 FILLER_4_711 ();
 sg13g2_decap_8 FILLER_4_718 ();
 sg13g2_decap_8 FILLER_4_725 ();
 sg13g2_decap_8 FILLER_4_732 ();
 sg13g2_decap_8 FILLER_4_739 ();
 sg13g2_decap_8 FILLER_4_746 ();
 sg13g2_decap_8 FILLER_4_753 ();
 sg13g2_decap_8 FILLER_4_760 ();
 sg13g2_decap_8 FILLER_4_767 ();
 sg13g2_decap_8 FILLER_4_774 ();
 sg13g2_decap_8 FILLER_4_781 ();
 sg13g2_decap_8 FILLER_4_788 ();
 sg13g2_decap_8 FILLER_4_795 ();
 sg13g2_decap_8 FILLER_4_802 ();
 sg13g2_decap_8 FILLER_4_809 ();
 sg13g2_decap_8 FILLER_4_816 ();
 sg13g2_decap_8 FILLER_4_823 ();
 sg13g2_decap_8 FILLER_4_830 ();
 sg13g2_decap_8 FILLER_4_837 ();
 sg13g2_decap_8 FILLER_4_844 ();
 sg13g2_decap_8 FILLER_4_851 ();
 sg13g2_decap_8 FILLER_4_858 ();
 sg13g2_decap_8 FILLER_4_865 ();
 sg13g2_decap_8 FILLER_4_872 ();
 sg13g2_decap_8 FILLER_4_879 ();
 sg13g2_decap_8 FILLER_4_886 ();
 sg13g2_decap_8 FILLER_4_893 ();
 sg13g2_decap_8 FILLER_4_900 ();
 sg13g2_decap_8 FILLER_4_907 ();
 sg13g2_decap_8 FILLER_4_914 ();
 sg13g2_decap_8 FILLER_4_921 ();
 sg13g2_decap_8 FILLER_4_928 ();
 sg13g2_decap_8 FILLER_4_935 ();
 sg13g2_decap_8 FILLER_4_942 ();
 sg13g2_decap_8 FILLER_4_949 ();
 sg13g2_decap_8 FILLER_4_956 ();
 sg13g2_decap_8 FILLER_4_963 ();
 sg13g2_decap_8 FILLER_4_970 ();
 sg13g2_decap_8 FILLER_4_977 ();
 sg13g2_decap_8 FILLER_4_984 ();
 sg13g2_decap_8 FILLER_4_991 ();
 sg13g2_decap_8 FILLER_4_998 ();
 sg13g2_decap_8 FILLER_4_1005 ();
 sg13g2_decap_8 FILLER_4_1012 ();
 sg13g2_decap_8 FILLER_4_1019 ();
 sg13g2_fill_2 FILLER_4_1026 ();
 sg13g2_fill_1 FILLER_4_1028 ();
 sg13g2_decap_8 FILLER_5_4 ();
 sg13g2_decap_8 FILLER_5_11 ();
 sg13g2_decap_8 FILLER_5_18 ();
 sg13g2_decap_8 FILLER_5_25 ();
 sg13g2_decap_8 FILLER_5_32 ();
 sg13g2_decap_8 FILLER_5_39 ();
 sg13g2_decap_8 FILLER_5_46 ();
 sg13g2_decap_8 FILLER_5_53 ();
 sg13g2_decap_8 FILLER_5_60 ();
 sg13g2_decap_8 FILLER_5_67 ();
 sg13g2_decap_8 FILLER_5_74 ();
 sg13g2_decap_8 FILLER_5_81 ();
 sg13g2_decap_8 FILLER_5_88 ();
 sg13g2_decap_8 FILLER_5_95 ();
 sg13g2_decap_8 FILLER_5_102 ();
 sg13g2_decap_8 FILLER_5_109 ();
 sg13g2_decap_8 FILLER_5_116 ();
 sg13g2_decap_8 FILLER_5_123 ();
 sg13g2_decap_8 FILLER_5_130 ();
 sg13g2_decap_8 FILLER_5_137 ();
 sg13g2_decap_8 FILLER_5_144 ();
 sg13g2_decap_8 FILLER_5_151 ();
 sg13g2_decap_8 FILLER_5_158 ();
 sg13g2_decap_8 FILLER_5_165 ();
 sg13g2_decap_8 FILLER_5_172 ();
 sg13g2_decap_8 FILLER_5_179 ();
 sg13g2_decap_8 FILLER_5_186 ();
 sg13g2_decap_8 FILLER_5_193 ();
 sg13g2_decap_8 FILLER_5_200 ();
 sg13g2_decap_8 FILLER_5_207 ();
 sg13g2_decap_8 FILLER_5_214 ();
 sg13g2_decap_8 FILLER_5_221 ();
 sg13g2_decap_8 FILLER_5_228 ();
 sg13g2_decap_8 FILLER_5_235 ();
 sg13g2_decap_8 FILLER_5_242 ();
 sg13g2_decap_8 FILLER_5_249 ();
 sg13g2_decap_8 FILLER_5_256 ();
 sg13g2_decap_8 FILLER_5_263 ();
 sg13g2_decap_8 FILLER_5_270 ();
 sg13g2_decap_8 FILLER_5_277 ();
 sg13g2_decap_8 FILLER_5_284 ();
 sg13g2_decap_8 FILLER_5_291 ();
 sg13g2_decap_8 FILLER_5_298 ();
 sg13g2_decap_8 FILLER_5_305 ();
 sg13g2_decap_8 FILLER_5_312 ();
 sg13g2_decap_8 FILLER_5_319 ();
 sg13g2_decap_8 FILLER_5_326 ();
 sg13g2_decap_8 FILLER_5_333 ();
 sg13g2_decap_8 FILLER_5_340 ();
 sg13g2_decap_8 FILLER_5_347 ();
 sg13g2_decap_8 FILLER_5_354 ();
 sg13g2_decap_8 FILLER_5_361 ();
 sg13g2_decap_8 FILLER_5_368 ();
 sg13g2_decap_8 FILLER_5_375 ();
 sg13g2_decap_8 FILLER_5_382 ();
 sg13g2_decap_8 FILLER_5_389 ();
 sg13g2_decap_8 FILLER_5_396 ();
 sg13g2_decap_8 FILLER_5_403 ();
 sg13g2_decap_8 FILLER_5_410 ();
 sg13g2_decap_8 FILLER_5_417 ();
 sg13g2_decap_8 FILLER_5_424 ();
 sg13g2_decap_8 FILLER_5_431 ();
 sg13g2_decap_8 FILLER_5_438 ();
 sg13g2_decap_8 FILLER_5_445 ();
 sg13g2_decap_8 FILLER_5_452 ();
 sg13g2_decap_8 FILLER_5_459 ();
 sg13g2_decap_8 FILLER_5_466 ();
 sg13g2_decap_8 FILLER_5_473 ();
 sg13g2_decap_8 FILLER_5_480 ();
 sg13g2_decap_8 FILLER_5_487 ();
 sg13g2_decap_8 FILLER_5_494 ();
 sg13g2_decap_8 FILLER_5_501 ();
 sg13g2_decap_8 FILLER_5_508 ();
 sg13g2_decap_8 FILLER_5_515 ();
 sg13g2_decap_8 FILLER_5_522 ();
 sg13g2_decap_8 FILLER_5_529 ();
 sg13g2_decap_8 FILLER_5_536 ();
 sg13g2_decap_8 FILLER_5_543 ();
 sg13g2_decap_8 FILLER_5_550 ();
 sg13g2_decap_8 FILLER_5_557 ();
 sg13g2_decap_8 FILLER_5_564 ();
 sg13g2_decap_8 FILLER_5_571 ();
 sg13g2_decap_8 FILLER_5_578 ();
 sg13g2_decap_8 FILLER_5_585 ();
 sg13g2_decap_8 FILLER_5_592 ();
 sg13g2_decap_8 FILLER_5_599 ();
 sg13g2_decap_8 FILLER_5_606 ();
 sg13g2_decap_8 FILLER_5_613 ();
 sg13g2_decap_8 FILLER_5_620 ();
 sg13g2_decap_8 FILLER_5_627 ();
 sg13g2_decap_8 FILLER_5_634 ();
 sg13g2_decap_8 FILLER_5_641 ();
 sg13g2_decap_8 FILLER_5_648 ();
 sg13g2_decap_8 FILLER_5_655 ();
 sg13g2_decap_8 FILLER_5_662 ();
 sg13g2_decap_8 FILLER_5_669 ();
 sg13g2_decap_8 FILLER_5_676 ();
 sg13g2_decap_8 FILLER_5_683 ();
 sg13g2_decap_8 FILLER_5_690 ();
 sg13g2_decap_8 FILLER_5_697 ();
 sg13g2_decap_8 FILLER_5_704 ();
 sg13g2_decap_8 FILLER_5_711 ();
 sg13g2_decap_8 FILLER_5_718 ();
 sg13g2_decap_8 FILLER_5_725 ();
 sg13g2_decap_8 FILLER_5_732 ();
 sg13g2_decap_8 FILLER_5_739 ();
 sg13g2_decap_8 FILLER_5_746 ();
 sg13g2_decap_8 FILLER_5_753 ();
 sg13g2_decap_8 FILLER_5_760 ();
 sg13g2_decap_8 FILLER_5_767 ();
 sg13g2_decap_8 FILLER_5_774 ();
 sg13g2_decap_8 FILLER_5_781 ();
 sg13g2_decap_8 FILLER_5_788 ();
 sg13g2_decap_8 FILLER_5_795 ();
 sg13g2_decap_8 FILLER_5_802 ();
 sg13g2_decap_8 FILLER_5_809 ();
 sg13g2_decap_8 FILLER_5_816 ();
 sg13g2_decap_8 FILLER_5_823 ();
 sg13g2_decap_8 FILLER_5_830 ();
 sg13g2_decap_8 FILLER_5_837 ();
 sg13g2_decap_8 FILLER_5_844 ();
 sg13g2_decap_8 FILLER_5_851 ();
 sg13g2_decap_8 FILLER_5_858 ();
 sg13g2_decap_8 FILLER_5_865 ();
 sg13g2_decap_8 FILLER_5_872 ();
 sg13g2_decap_8 FILLER_5_879 ();
 sg13g2_decap_8 FILLER_5_886 ();
 sg13g2_decap_8 FILLER_5_893 ();
 sg13g2_decap_8 FILLER_5_900 ();
 sg13g2_decap_8 FILLER_5_907 ();
 sg13g2_decap_8 FILLER_5_914 ();
 sg13g2_decap_8 FILLER_5_921 ();
 sg13g2_decap_8 FILLER_5_928 ();
 sg13g2_decap_8 FILLER_5_935 ();
 sg13g2_decap_8 FILLER_5_942 ();
 sg13g2_decap_8 FILLER_5_949 ();
 sg13g2_decap_8 FILLER_5_956 ();
 sg13g2_decap_8 FILLER_5_963 ();
 sg13g2_decap_8 FILLER_5_970 ();
 sg13g2_decap_8 FILLER_5_977 ();
 sg13g2_decap_8 FILLER_5_984 ();
 sg13g2_decap_8 FILLER_5_991 ();
 sg13g2_decap_8 FILLER_5_998 ();
 sg13g2_decap_8 FILLER_5_1005 ();
 sg13g2_decap_8 FILLER_5_1012 ();
 sg13g2_decap_8 FILLER_5_1019 ();
 sg13g2_fill_2 FILLER_5_1026 ();
 sg13g2_fill_1 FILLER_5_1028 ();
 sg13g2_decap_8 FILLER_6_4 ();
 sg13g2_decap_8 FILLER_6_11 ();
 sg13g2_decap_8 FILLER_6_18 ();
 sg13g2_decap_8 FILLER_6_25 ();
 sg13g2_decap_8 FILLER_6_32 ();
 sg13g2_decap_8 FILLER_6_39 ();
 sg13g2_decap_8 FILLER_6_46 ();
 sg13g2_decap_8 FILLER_6_53 ();
 sg13g2_decap_8 FILLER_6_60 ();
 sg13g2_decap_8 FILLER_6_67 ();
 sg13g2_decap_8 FILLER_6_74 ();
 sg13g2_decap_8 FILLER_6_81 ();
 sg13g2_decap_8 FILLER_6_88 ();
 sg13g2_decap_8 FILLER_6_95 ();
 sg13g2_decap_8 FILLER_6_102 ();
 sg13g2_decap_8 FILLER_6_109 ();
 sg13g2_decap_8 FILLER_6_116 ();
 sg13g2_decap_8 FILLER_6_123 ();
 sg13g2_decap_8 FILLER_6_130 ();
 sg13g2_decap_8 FILLER_6_137 ();
 sg13g2_decap_8 FILLER_6_144 ();
 sg13g2_decap_8 FILLER_6_151 ();
 sg13g2_decap_8 FILLER_6_158 ();
 sg13g2_decap_8 FILLER_6_165 ();
 sg13g2_decap_8 FILLER_6_172 ();
 sg13g2_decap_8 FILLER_6_179 ();
 sg13g2_decap_8 FILLER_6_186 ();
 sg13g2_decap_8 FILLER_6_193 ();
 sg13g2_decap_8 FILLER_6_200 ();
 sg13g2_decap_8 FILLER_6_207 ();
 sg13g2_decap_8 FILLER_6_214 ();
 sg13g2_decap_8 FILLER_6_221 ();
 sg13g2_decap_8 FILLER_6_228 ();
 sg13g2_decap_8 FILLER_6_235 ();
 sg13g2_decap_8 FILLER_6_242 ();
 sg13g2_decap_8 FILLER_6_249 ();
 sg13g2_decap_8 FILLER_6_256 ();
 sg13g2_decap_8 FILLER_6_263 ();
 sg13g2_decap_8 FILLER_6_270 ();
 sg13g2_decap_8 FILLER_6_277 ();
 sg13g2_decap_8 FILLER_6_284 ();
 sg13g2_decap_8 FILLER_6_291 ();
 sg13g2_decap_8 FILLER_6_298 ();
 sg13g2_decap_8 FILLER_6_305 ();
 sg13g2_decap_8 FILLER_6_312 ();
 sg13g2_decap_8 FILLER_6_319 ();
 sg13g2_decap_8 FILLER_6_326 ();
 sg13g2_decap_8 FILLER_6_333 ();
 sg13g2_decap_8 FILLER_6_340 ();
 sg13g2_decap_8 FILLER_6_347 ();
 sg13g2_decap_8 FILLER_6_354 ();
 sg13g2_decap_8 FILLER_6_361 ();
 sg13g2_decap_8 FILLER_6_368 ();
 sg13g2_decap_8 FILLER_6_375 ();
 sg13g2_decap_8 FILLER_6_382 ();
 sg13g2_decap_8 FILLER_6_389 ();
 sg13g2_decap_8 FILLER_6_396 ();
 sg13g2_decap_8 FILLER_6_403 ();
 sg13g2_decap_8 FILLER_6_410 ();
 sg13g2_decap_8 FILLER_6_417 ();
 sg13g2_decap_8 FILLER_6_424 ();
 sg13g2_decap_8 FILLER_6_431 ();
 sg13g2_decap_8 FILLER_6_438 ();
 sg13g2_decap_8 FILLER_6_445 ();
 sg13g2_decap_8 FILLER_6_452 ();
 sg13g2_decap_8 FILLER_6_459 ();
 sg13g2_decap_8 FILLER_6_466 ();
 sg13g2_decap_8 FILLER_6_473 ();
 sg13g2_decap_8 FILLER_6_480 ();
 sg13g2_decap_8 FILLER_6_487 ();
 sg13g2_decap_8 FILLER_6_494 ();
 sg13g2_decap_8 FILLER_6_501 ();
 sg13g2_decap_8 FILLER_6_508 ();
 sg13g2_decap_8 FILLER_6_515 ();
 sg13g2_decap_8 FILLER_6_522 ();
 sg13g2_decap_8 FILLER_6_529 ();
 sg13g2_decap_8 FILLER_6_536 ();
 sg13g2_decap_8 FILLER_6_543 ();
 sg13g2_decap_8 FILLER_6_550 ();
 sg13g2_decap_8 FILLER_6_557 ();
 sg13g2_decap_8 FILLER_6_564 ();
 sg13g2_decap_8 FILLER_6_571 ();
 sg13g2_decap_8 FILLER_6_578 ();
 sg13g2_decap_8 FILLER_6_585 ();
 sg13g2_decap_8 FILLER_6_592 ();
 sg13g2_decap_8 FILLER_6_599 ();
 sg13g2_decap_8 FILLER_6_606 ();
 sg13g2_decap_8 FILLER_6_613 ();
 sg13g2_decap_8 FILLER_6_620 ();
 sg13g2_decap_8 FILLER_6_627 ();
 sg13g2_decap_8 FILLER_6_634 ();
 sg13g2_decap_8 FILLER_6_641 ();
 sg13g2_decap_8 FILLER_6_648 ();
 sg13g2_decap_8 FILLER_6_655 ();
 sg13g2_decap_8 FILLER_6_662 ();
 sg13g2_decap_8 FILLER_6_669 ();
 sg13g2_decap_8 FILLER_6_676 ();
 sg13g2_decap_8 FILLER_6_683 ();
 sg13g2_decap_8 FILLER_6_690 ();
 sg13g2_decap_8 FILLER_6_697 ();
 sg13g2_decap_8 FILLER_6_704 ();
 sg13g2_decap_8 FILLER_6_711 ();
 sg13g2_decap_8 FILLER_6_718 ();
 sg13g2_decap_8 FILLER_6_725 ();
 sg13g2_decap_8 FILLER_6_732 ();
 sg13g2_decap_8 FILLER_6_739 ();
 sg13g2_decap_8 FILLER_6_746 ();
 sg13g2_decap_8 FILLER_6_753 ();
 sg13g2_decap_8 FILLER_6_760 ();
 sg13g2_decap_8 FILLER_6_767 ();
 sg13g2_decap_8 FILLER_6_774 ();
 sg13g2_decap_8 FILLER_6_781 ();
 sg13g2_decap_8 FILLER_6_788 ();
 sg13g2_decap_8 FILLER_6_795 ();
 sg13g2_decap_8 FILLER_6_802 ();
 sg13g2_decap_8 FILLER_6_809 ();
 sg13g2_decap_8 FILLER_6_816 ();
 sg13g2_decap_8 FILLER_6_823 ();
 sg13g2_decap_8 FILLER_6_830 ();
 sg13g2_decap_8 FILLER_6_837 ();
 sg13g2_decap_8 FILLER_6_844 ();
 sg13g2_decap_8 FILLER_6_851 ();
 sg13g2_decap_8 FILLER_6_858 ();
 sg13g2_decap_8 FILLER_6_865 ();
 sg13g2_decap_8 FILLER_6_872 ();
 sg13g2_decap_8 FILLER_6_879 ();
 sg13g2_decap_8 FILLER_6_886 ();
 sg13g2_decap_8 FILLER_6_893 ();
 sg13g2_decap_8 FILLER_6_900 ();
 sg13g2_decap_8 FILLER_6_907 ();
 sg13g2_decap_8 FILLER_6_914 ();
 sg13g2_decap_8 FILLER_6_921 ();
 sg13g2_decap_8 FILLER_6_928 ();
 sg13g2_decap_8 FILLER_6_935 ();
 sg13g2_decap_8 FILLER_6_942 ();
 sg13g2_decap_8 FILLER_6_949 ();
 sg13g2_decap_8 FILLER_6_956 ();
 sg13g2_decap_8 FILLER_6_963 ();
 sg13g2_decap_8 FILLER_6_970 ();
 sg13g2_decap_8 FILLER_6_977 ();
 sg13g2_decap_8 FILLER_6_984 ();
 sg13g2_decap_8 FILLER_6_991 ();
 sg13g2_decap_8 FILLER_6_998 ();
 sg13g2_decap_8 FILLER_6_1005 ();
 sg13g2_decap_8 FILLER_6_1012 ();
 sg13g2_decap_8 FILLER_6_1019 ();
 sg13g2_fill_2 FILLER_6_1026 ();
 sg13g2_fill_1 FILLER_6_1028 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_decap_8 FILLER_7_406 ();
 sg13g2_decap_8 FILLER_7_413 ();
 sg13g2_decap_8 FILLER_7_420 ();
 sg13g2_decap_8 FILLER_7_427 ();
 sg13g2_decap_8 FILLER_7_434 ();
 sg13g2_decap_8 FILLER_7_441 ();
 sg13g2_decap_8 FILLER_7_448 ();
 sg13g2_decap_8 FILLER_7_455 ();
 sg13g2_decap_8 FILLER_7_462 ();
 sg13g2_decap_8 FILLER_7_469 ();
 sg13g2_decap_8 FILLER_7_476 ();
 sg13g2_decap_8 FILLER_7_483 ();
 sg13g2_decap_8 FILLER_7_490 ();
 sg13g2_decap_8 FILLER_7_497 ();
 sg13g2_decap_8 FILLER_7_504 ();
 sg13g2_decap_8 FILLER_7_511 ();
 sg13g2_decap_8 FILLER_7_518 ();
 sg13g2_decap_8 FILLER_7_525 ();
 sg13g2_decap_8 FILLER_7_532 ();
 sg13g2_decap_8 FILLER_7_539 ();
 sg13g2_decap_8 FILLER_7_546 ();
 sg13g2_decap_8 FILLER_7_553 ();
 sg13g2_decap_8 FILLER_7_560 ();
 sg13g2_decap_8 FILLER_7_567 ();
 sg13g2_decap_8 FILLER_7_574 ();
 sg13g2_decap_8 FILLER_7_581 ();
 sg13g2_decap_8 FILLER_7_588 ();
 sg13g2_decap_8 FILLER_7_595 ();
 sg13g2_decap_8 FILLER_7_602 ();
 sg13g2_decap_8 FILLER_7_609 ();
 sg13g2_decap_8 FILLER_7_616 ();
 sg13g2_decap_8 FILLER_7_623 ();
 sg13g2_decap_8 FILLER_7_630 ();
 sg13g2_decap_8 FILLER_7_637 ();
 sg13g2_decap_8 FILLER_7_644 ();
 sg13g2_decap_8 FILLER_7_651 ();
 sg13g2_decap_8 FILLER_7_658 ();
 sg13g2_decap_8 FILLER_7_665 ();
 sg13g2_decap_8 FILLER_7_672 ();
 sg13g2_decap_8 FILLER_7_679 ();
 sg13g2_decap_8 FILLER_7_686 ();
 sg13g2_decap_8 FILLER_7_693 ();
 sg13g2_decap_8 FILLER_7_700 ();
 sg13g2_decap_8 FILLER_7_707 ();
 sg13g2_decap_8 FILLER_7_714 ();
 sg13g2_decap_8 FILLER_7_721 ();
 sg13g2_decap_8 FILLER_7_728 ();
 sg13g2_decap_8 FILLER_7_735 ();
 sg13g2_decap_8 FILLER_7_742 ();
 sg13g2_decap_8 FILLER_7_749 ();
 sg13g2_decap_8 FILLER_7_756 ();
 sg13g2_decap_8 FILLER_7_763 ();
 sg13g2_decap_8 FILLER_7_770 ();
 sg13g2_decap_8 FILLER_7_777 ();
 sg13g2_decap_8 FILLER_7_784 ();
 sg13g2_decap_8 FILLER_7_791 ();
 sg13g2_decap_8 FILLER_7_798 ();
 sg13g2_decap_8 FILLER_7_805 ();
 sg13g2_decap_8 FILLER_7_812 ();
 sg13g2_decap_8 FILLER_7_819 ();
 sg13g2_decap_8 FILLER_7_826 ();
 sg13g2_decap_8 FILLER_7_833 ();
 sg13g2_decap_8 FILLER_7_840 ();
 sg13g2_decap_8 FILLER_7_847 ();
 sg13g2_decap_8 FILLER_7_854 ();
 sg13g2_decap_8 FILLER_7_861 ();
 sg13g2_decap_8 FILLER_7_868 ();
 sg13g2_decap_8 FILLER_7_875 ();
 sg13g2_decap_8 FILLER_7_882 ();
 sg13g2_decap_8 FILLER_7_889 ();
 sg13g2_decap_8 FILLER_7_896 ();
 sg13g2_decap_8 FILLER_7_903 ();
 sg13g2_decap_8 FILLER_7_910 ();
 sg13g2_decap_8 FILLER_7_917 ();
 sg13g2_decap_8 FILLER_7_924 ();
 sg13g2_decap_8 FILLER_7_931 ();
 sg13g2_decap_8 FILLER_7_938 ();
 sg13g2_decap_8 FILLER_7_945 ();
 sg13g2_decap_8 FILLER_7_952 ();
 sg13g2_decap_8 FILLER_7_959 ();
 sg13g2_decap_8 FILLER_7_966 ();
 sg13g2_decap_8 FILLER_7_973 ();
 sg13g2_decap_8 FILLER_7_980 ();
 sg13g2_decap_8 FILLER_7_987 ();
 sg13g2_decap_8 FILLER_7_994 ();
 sg13g2_decap_8 FILLER_7_1001 ();
 sg13g2_decap_8 FILLER_7_1008 ();
 sg13g2_decap_8 FILLER_7_1015 ();
 sg13g2_decap_8 FILLER_7_1022 ();
 sg13g2_decap_8 FILLER_8_4 ();
 sg13g2_decap_8 FILLER_8_11 ();
 sg13g2_decap_8 FILLER_8_18 ();
 sg13g2_decap_8 FILLER_8_25 ();
 sg13g2_decap_8 FILLER_8_32 ();
 sg13g2_decap_8 FILLER_8_39 ();
 sg13g2_decap_8 FILLER_8_46 ();
 sg13g2_decap_8 FILLER_8_53 ();
 sg13g2_decap_8 FILLER_8_60 ();
 sg13g2_decap_8 FILLER_8_67 ();
 sg13g2_decap_8 FILLER_8_74 ();
 sg13g2_decap_8 FILLER_8_81 ();
 sg13g2_decap_8 FILLER_8_88 ();
 sg13g2_decap_8 FILLER_8_95 ();
 sg13g2_decap_8 FILLER_8_102 ();
 sg13g2_decap_8 FILLER_8_109 ();
 sg13g2_decap_8 FILLER_8_116 ();
 sg13g2_decap_8 FILLER_8_123 ();
 sg13g2_decap_8 FILLER_8_130 ();
 sg13g2_decap_8 FILLER_8_137 ();
 sg13g2_decap_8 FILLER_8_144 ();
 sg13g2_decap_8 FILLER_8_151 ();
 sg13g2_decap_8 FILLER_8_158 ();
 sg13g2_decap_8 FILLER_8_165 ();
 sg13g2_decap_8 FILLER_8_172 ();
 sg13g2_decap_8 FILLER_8_179 ();
 sg13g2_decap_8 FILLER_8_186 ();
 sg13g2_decap_8 FILLER_8_193 ();
 sg13g2_decap_8 FILLER_8_200 ();
 sg13g2_decap_8 FILLER_8_207 ();
 sg13g2_decap_8 FILLER_8_214 ();
 sg13g2_decap_8 FILLER_8_221 ();
 sg13g2_decap_8 FILLER_8_228 ();
 sg13g2_decap_8 FILLER_8_235 ();
 sg13g2_decap_8 FILLER_8_242 ();
 sg13g2_decap_8 FILLER_8_249 ();
 sg13g2_decap_8 FILLER_8_256 ();
 sg13g2_decap_8 FILLER_8_263 ();
 sg13g2_decap_8 FILLER_8_270 ();
 sg13g2_decap_8 FILLER_8_277 ();
 sg13g2_decap_8 FILLER_8_284 ();
 sg13g2_decap_8 FILLER_8_291 ();
 sg13g2_decap_8 FILLER_8_298 ();
 sg13g2_decap_8 FILLER_8_305 ();
 sg13g2_decap_8 FILLER_8_312 ();
 sg13g2_decap_8 FILLER_8_319 ();
 sg13g2_decap_8 FILLER_8_326 ();
 sg13g2_decap_8 FILLER_8_333 ();
 sg13g2_decap_8 FILLER_8_340 ();
 sg13g2_decap_8 FILLER_8_347 ();
 sg13g2_decap_8 FILLER_8_354 ();
 sg13g2_decap_8 FILLER_8_361 ();
 sg13g2_decap_8 FILLER_8_368 ();
 sg13g2_decap_8 FILLER_8_375 ();
 sg13g2_decap_8 FILLER_8_382 ();
 sg13g2_decap_8 FILLER_8_389 ();
 sg13g2_decap_8 FILLER_8_396 ();
 sg13g2_decap_8 FILLER_8_403 ();
 sg13g2_decap_8 FILLER_8_410 ();
 sg13g2_decap_8 FILLER_8_417 ();
 sg13g2_decap_8 FILLER_8_424 ();
 sg13g2_decap_8 FILLER_8_431 ();
 sg13g2_decap_8 FILLER_8_438 ();
 sg13g2_decap_8 FILLER_8_445 ();
 sg13g2_decap_8 FILLER_8_452 ();
 sg13g2_decap_8 FILLER_8_459 ();
 sg13g2_decap_8 FILLER_8_466 ();
 sg13g2_decap_8 FILLER_8_473 ();
 sg13g2_decap_8 FILLER_8_480 ();
 sg13g2_decap_8 FILLER_8_487 ();
 sg13g2_decap_8 FILLER_8_494 ();
 sg13g2_decap_8 FILLER_8_501 ();
 sg13g2_decap_8 FILLER_8_508 ();
 sg13g2_decap_8 FILLER_8_515 ();
 sg13g2_decap_8 FILLER_8_522 ();
 sg13g2_decap_8 FILLER_8_529 ();
 sg13g2_decap_8 FILLER_8_536 ();
 sg13g2_decap_8 FILLER_8_543 ();
 sg13g2_decap_8 FILLER_8_550 ();
 sg13g2_decap_8 FILLER_8_557 ();
 sg13g2_decap_8 FILLER_8_564 ();
 sg13g2_decap_8 FILLER_8_571 ();
 sg13g2_decap_8 FILLER_8_578 ();
 sg13g2_decap_8 FILLER_8_585 ();
 sg13g2_decap_8 FILLER_8_592 ();
 sg13g2_decap_8 FILLER_8_599 ();
 sg13g2_decap_8 FILLER_8_606 ();
 sg13g2_decap_8 FILLER_8_613 ();
 sg13g2_decap_8 FILLER_8_620 ();
 sg13g2_decap_8 FILLER_8_627 ();
 sg13g2_decap_8 FILLER_8_634 ();
 sg13g2_decap_8 FILLER_8_641 ();
 sg13g2_decap_8 FILLER_8_648 ();
 sg13g2_decap_8 FILLER_8_655 ();
 sg13g2_decap_8 FILLER_8_662 ();
 sg13g2_decap_8 FILLER_8_669 ();
 sg13g2_decap_8 FILLER_8_676 ();
 sg13g2_decap_8 FILLER_8_683 ();
 sg13g2_decap_8 FILLER_8_690 ();
 sg13g2_decap_8 FILLER_8_697 ();
 sg13g2_decap_8 FILLER_8_704 ();
 sg13g2_decap_8 FILLER_8_711 ();
 sg13g2_decap_8 FILLER_8_718 ();
 sg13g2_decap_8 FILLER_8_725 ();
 sg13g2_decap_8 FILLER_8_732 ();
 sg13g2_decap_8 FILLER_8_739 ();
 sg13g2_decap_8 FILLER_8_746 ();
 sg13g2_decap_8 FILLER_8_753 ();
 sg13g2_decap_8 FILLER_8_760 ();
 sg13g2_decap_8 FILLER_8_767 ();
 sg13g2_decap_8 FILLER_8_774 ();
 sg13g2_decap_8 FILLER_8_781 ();
 sg13g2_decap_8 FILLER_8_788 ();
 sg13g2_decap_8 FILLER_8_795 ();
 sg13g2_decap_8 FILLER_8_802 ();
 sg13g2_decap_8 FILLER_8_809 ();
 sg13g2_decap_8 FILLER_8_816 ();
 sg13g2_decap_8 FILLER_8_823 ();
 sg13g2_decap_8 FILLER_8_830 ();
 sg13g2_decap_8 FILLER_8_837 ();
 sg13g2_decap_8 FILLER_8_844 ();
 sg13g2_decap_8 FILLER_8_851 ();
 sg13g2_decap_8 FILLER_8_858 ();
 sg13g2_decap_8 FILLER_8_865 ();
 sg13g2_decap_8 FILLER_8_872 ();
 sg13g2_decap_8 FILLER_8_879 ();
 sg13g2_decap_8 FILLER_8_886 ();
 sg13g2_decap_8 FILLER_8_893 ();
 sg13g2_decap_8 FILLER_8_900 ();
 sg13g2_decap_8 FILLER_8_907 ();
 sg13g2_decap_8 FILLER_8_914 ();
 sg13g2_decap_8 FILLER_8_921 ();
 sg13g2_decap_8 FILLER_8_928 ();
 sg13g2_decap_8 FILLER_8_935 ();
 sg13g2_decap_8 FILLER_8_942 ();
 sg13g2_decap_8 FILLER_8_949 ();
 sg13g2_decap_8 FILLER_8_956 ();
 sg13g2_decap_8 FILLER_8_963 ();
 sg13g2_decap_8 FILLER_8_970 ();
 sg13g2_decap_8 FILLER_8_977 ();
 sg13g2_decap_8 FILLER_8_984 ();
 sg13g2_decap_8 FILLER_8_991 ();
 sg13g2_decap_8 FILLER_8_998 ();
 sg13g2_decap_8 FILLER_8_1005 ();
 sg13g2_decap_8 FILLER_8_1012 ();
 sg13g2_decap_8 FILLER_8_1019 ();
 sg13g2_fill_2 FILLER_8_1026 ();
 sg13g2_fill_1 FILLER_8_1028 ();
 sg13g2_decap_8 FILLER_9_4 ();
 sg13g2_decap_8 FILLER_9_11 ();
 sg13g2_decap_8 FILLER_9_18 ();
 sg13g2_decap_8 FILLER_9_25 ();
 sg13g2_decap_8 FILLER_9_32 ();
 sg13g2_decap_8 FILLER_9_39 ();
 sg13g2_decap_8 FILLER_9_46 ();
 sg13g2_decap_8 FILLER_9_53 ();
 sg13g2_decap_8 FILLER_9_60 ();
 sg13g2_decap_8 FILLER_9_67 ();
 sg13g2_decap_8 FILLER_9_74 ();
 sg13g2_decap_8 FILLER_9_81 ();
 sg13g2_decap_8 FILLER_9_88 ();
 sg13g2_decap_8 FILLER_9_95 ();
 sg13g2_decap_8 FILLER_9_102 ();
 sg13g2_decap_8 FILLER_9_109 ();
 sg13g2_decap_8 FILLER_9_116 ();
 sg13g2_decap_8 FILLER_9_123 ();
 sg13g2_decap_8 FILLER_9_130 ();
 sg13g2_decap_8 FILLER_9_137 ();
 sg13g2_decap_8 FILLER_9_144 ();
 sg13g2_decap_8 FILLER_9_151 ();
 sg13g2_decap_8 FILLER_9_158 ();
 sg13g2_decap_8 FILLER_9_165 ();
 sg13g2_decap_8 FILLER_9_172 ();
 sg13g2_decap_8 FILLER_9_179 ();
 sg13g2_decap_8 FILLER_9_186 ();
 sg13g2_decap_8 FILLER_9_193 ();
 sg13g2_decap_8 FILLER_9_200 ();
 sg13g2_decap_8 FILLER_9_207 ();
 sg13g2_decap_8 FILLER_9_214 ();
 sg13g2_decap_8 FILLER_9_221 ();
 sg13g2_decap_8 FILLER_9_228 ();
 sg13g2_decap_8 FILLER_9_235 ();
 sg13g2_decap_8 FILLER_9_242 ();
 sg13g2_decap_8 FILLER_9_249 ();
 sg13g2_decap_8 FILLER_9_256 ();
 sg13g2_decap_8 FILLER_9_263 ();
 sg13g2_decap_8 FILLER_9_270 ();
 sg13g2_decap_8 FILLER_9_277 ();
 sg13g2_decap_8 FILLER_9_284 ();
 sg13g2_decap_8 FILLER_9_291 ();
 sg13g2_decap_8 FILLER_9_298 ();
 sg13g2_decap_8 FILLER_9_305 ();
 sg13g2_decap_8 FILLER_9_312 ();
 sg13g2_decap_8 FILLER_9_319 ();
 sg13g2_decap_8 FILLER_9_326 ();
 sg13g2_decap_8 FILLER_9_333 ();
 sg13g2_decap_8 FILLER_9_340 ();
 sg13g2_decap_8 FILLER_9_347 ();
 sg13g2_decap_8 FILLER_9_354 ();
 sg13g2_decap_8 FILLER_9_361 ();
 sg13g2_decap_8 FILLER_9_368 ();
 sg13g2_decap_8 FILLER_9_375 ();
 sg13g2_decap_8 FILLER_9_382 ();
 sg13g2_decap_8 FILLER_9_389 ();
 sg13g2_decap_8 FILLER_9_396 ();
 sg13g2_decap_8 FILLER_9_403 ();
 sg13g2_decap_8 FILLER_9_410 ();
 sg13g2_decap_8 FILLER_9_417 ();
 sg13g2_decap_8 FILLER_9_424 ();
 sg13g2_decap_8 FILLER_9_431 ();
 sg13g2_decap_8 FILLER_9_438 ();
 sg13g2_decap_8 FILLER_9_445 ();
 sg13g2_decap_8 FILLER_9_452 ();
 sg13g2_decap_8 FILLER_9_459 ();
 sg13g2_decap_8 FILLER_9_466 ();
 sg13g2_decap_8 FILLER_9_473 ();
 sg13g2_decap_8 FILLER_9_480 ();
 sg13g2_decap_8 FILLER_9_487 ();
 sg13g2_decap_8 FILLER_9_494 ();
 sg13g2_decap_8 FILLER_9_501 ();
 sg13g2_decap_8 FILLER_9_508 ();
 sg13g2_decap_8 FILLER_9_515 ();
 sg13g2_decap_8 FILLER_9_522 ();
 sg13g2_decap_8 FILLER_9_529 ();
 sg13g2_decap_8 FILLER_9_536 ();
 sg13g2_decap_8 FILLER_9_543 ();
 sg13g2_decap_8 FILLER_9_550 ();
 sg13g2_decap_8 FILLER_9_557 ();
 sg13g2_decap_8 FILLER_9_564 ();
 sg13g2_decap_8 FILLER_9_571 ();
 sg13g2_decap_8 FILLER_9_578 ();
 sg13g2_decap_8 FILLER_9_585 ();
 sg13g2_decap_8 FILLER_9_592 ();
 sg13g2_decap_8 FILLER_9_599 ();
 sg13g2_decap_8 FILLER_9_606 ();
 sg13g2_decap_8 FILLER_9_613 ();
 sg13g2_decap_8 FILLER_9_620 ();
 sg13g2_decap_8 FILLER_9_627 ();
 sg13g2_decap_8 FILLER_9_634 ();
 sg13g2_decap_8 FILLER_9_641 ();
 sg13g2_decap_8 FILLER_9_648 ();
 sg13g2_decap_8 FILLER_9_655 ();
 sg13g2_decap_8 FILLER_9_662 ();
 sg13g2_decap_8 FILLER_9_669 ();
 sg13g2_decap_8 FILLER_9_676 ();
 sg13g2_decap_8 FILLER_9_683 ();
 sg13g2_decap_8 FILLER_9_690 ();
 sg13g2_decap_8 FILLER_9_697 ();
 sg13g2_decap_8 FILLER_9_704 ();
 sg13g2_decap_8 FILLER_9_711 ();
 sg13g2_decap_8 FILLER_9_718 ();
 sg13g2_decap_8 FILLER_9_725 ();
 sg13g2_decap_8 FILLER_9_732 ();
 sg13g2_decap_8 FILLER_9_739 ();
 sg13g2_decap_8 FILLER_9_746 ();
 sg13g2_decap_8 FILLER_9_753 ();
 sg13g2_decap_8 FILLER_9_760 ();
 sg13g2_decap_8 FILLER_9_767 ();
 sg13g2_decap_8 FILLER_9_774 ();
 sg13g2_decap_8 FILLER_9_781 ();
 sg13g2_decap_8 FILLER_9_788 ();
 sg13g2_decap_8 FILLER_9_795 ();
 sg13g2_decap_8 FILLER_9_802 ();
 sg13g2_decap_8 FILLER_9_809 ();
 sg13g2_decap_8 FILLER_9_816 ();
 sg13g2_decap_8 FILLER_9_823 ();
 sg13g2_decap_8 FILLER_9_830 ();
 sg13g2_decap_8 FILLER_9_837 ();
 sg13g2_decap_8 FILLER_9_844 ();
 sg13g2_decap_8 FILLER_9_851 ();
 sg13g2_decap_8 FILLER_9_858 ();
 sg13g2_decap_8 FILLER_9_865 ();
 sg13g2_decap_8 FILLER_9_872 ();
 sg13g2_decap_8 FILLER_9_879 ();
 sg13g2_decap_8 FILLER_9_886 ();
 sg13g2_decap_8 FILLER_9_893 ();
 sg13g2_decap_8 FILLER_9_900 ();
 sg13g2_decap_8 FILLER_9_907 ();
 sg13g2_decap_8 FILLER_9_914 ();
 sg13g2_decap_8 FILLER_9_921 ();
 sg13g2_decap_8 FILLER_9_928 ();
 sg13g2_decap_8 FILLER_9_935 ();
 sg13g2_decap_8 FILLER_9_942 ();
 sg13g2_decap_8 FILLER_9_949 ();
 sg13g2_decap_8 FILLER_9_956 ();
 sg13g2_decap_8 FILLER_9_963 ();
 sg13g2_decap_8 FILLER_9_970 ();
 sg13g2_decap_8 FILLER_9_977 ();
 sg13g2_decap_8 FILLER_9_984 ();
 sg13g2_decap_8 FILLER_9_991 ();
 sg13g2_decap_8 FILLER_9_998 ();
 sg13g2_decap_8 FILLER_9_1005 ();
 sg13g2_decap_8 FILLER_9_1012 ();
 sg13g2_decap_8 FILLER_9_1019 ();
 sg13g2_fill_2 FILLER_9_1026 ();
 sg13g2_fill_1 FILLER_9_1028 ();
 sg13g2_decap_8 FILLER_10_4 ();
 sg13g2_decap_8 FILLER_10_11 ();
 sg13g2_decap_8 FILLER_10_18 ();
 sg13g2_decap_8 FILLER_10_25 ();
 sg13g2_decap_8 FILLER_10_32 ();
 sg13g2_decap_8 FILLER_10_39 ();
 sg13g2_decap_8 FILLER_10_46 ();
 sg13g2_decap_8 FILLER_10_53 ();
 sg13g2_decap_8 FILLER_10_60 ();
 sg13g2_decap_8 FILLER_10_67 ();
 sg13g2_decap_8 FILLER_10_74 ();
 sg13g2_decap_8 FILLER_10_81 ();
 sg13g2_decap_8 FILLER_10_88 ();
 sg13g2_decap_8 FILLER_10_95 ();
 sg13g2_decap_8 FILLER_10_102 ();
 sg13g2_decap_8 FILLER_10_109 ();
 sg13g2_decap_8 FILLER_10_116 ();
 sg13g2_decap_8 FILLER_10_123 ();
 sg13g2_decap_8 FILLER_10_130 ();
 sg13g2_decap_8 FILLER_10_137 ();
 sg13g2_decap_8 FILLER_10_144 ();
 sg13g2_decap_8 FILLER_10_151 ();
 sg13g2_decap_8 FILLER_10_158 ();
 sg13g2_decap_8 FILLER_10_165 ();
 sg13g2_decap_8 FILLER_10_172 ();
 sg13g2_decap_8 FILLER_10_179 ();
 sg13g2_decap_8 FILLER_10_186 ();
 sg13g2_decap_8 FILLER_10_193 ();
 sg13g2_decap_8 FILLER_10_200 ();
 sg13g2_decap_8 FILLER_10_207 ();
 sg13g2_decap_8 FILLER_10_214 ();
 sg13g2_decap_8 FILLER_10_221 ();
 sg13g2_decap_8 FILLER_10_228 ();
 sg13g2_decap_8 FILLER_10_235 ();
 sg13g2_decap_8 FILLER_10_242 ();
 sg13g2_decap_8 FILLER_10_249 ();
 sg13g2_decap_8 FILLER_10_256 ();
 sg13g2_decap_8 FILLER_10_263 ();
 sg13g2_decap_8 FILLER_10_270 ();
 sg13g2_decap_8 FILLER_10_277 ();
 sg13g2_decap_8 FILLER_10_284 ();
 sg13g2_decap_8 FILLER_10_291 ();
 sg13g2_decap_8 FILLER_10_298 ();
 sg13g2_decap_8 FILLER_10_305 ();
 sg13g2_decap_8 FILLER_10_312 ();
 sg13g2_decap_8 FILLER_10_319 ();
 sg13g2_decap_8 FILLER_10_326 ();
 sg13g2_decap_8 FILLER_10_333 ();
 sg13g2_decap_8 FILLER_10_340 ();
 sg13g2_decap_8 FILLER_10_347 ();
 sg13g2_decap_8 FILLER_10_354 ();
 sg13g2_decap_8 FILLER_10_361 ();
 sg13g2_decap_8 FILLER_10_368 ();
 sg13g2_decap_8 FILLER_10_375 ();
 sg13g2_decap_8 FILLER_10_382 ();
 sg13g2_decap_8 FILLER_10_389 ();
 sg13g2_decap_8 FILLER_10_396 ();
 sg13g2_decap_8 FILLER_10_403 ();
 sg13g2_decap_8 FILLER_10_410 ();
 sg13g2_decap_8 FILLER_10_417 ();
 sg13g2_decap_8 FILLER_10_424 ();
 sg13g2_decap_8 FILLER_10_431 ();
 sg13g2_decap_8 FILLER_10_438 ();
 sg13g2_decap_8 FILLER_10_445 ();
 sg13g2_decap_8 FILLER_10_452 ();
 sg13g2_decap_8 FILLER_10_459 ();
 sg13g2_decap_8 FILLER_10_466 ();
 sg13g2_decap_8 FILLER_10_473 ();
 sg13g2_decap_8 FILLER_10_480 ();
 sg13g2_decap_8 FILLER_10_487 ();
 sg13g2_decap_8 FILLER_10_494 ();
 sg13g2_decap_8 FILLER_10_501 ();
 sg13g2_decap_8 FILLER_10_508 ();
 sg13g2_decap_8 FILLER_10_515 ();
 sg13g2_decap_8 FILLER_10_522 ();
 sg13g2_decap_8 FILLER_10_529 ();
 sg13g2_decap_8 FILLER_10_536 ();
 sg13g2_decap_8 FILLER_10_543 ();
 sg13g2_decap_8 FILLER_10_550 ();
 sg13g2_decap_8 FILLER_10_557 ();
 sg13g2_decap_8 FILLER_10_564 ();
 sg13g2_decap_8 FILLER_10_571 ();
 sg13g2_decap_8 FILLER_10_578 ();
 sg13g2_decap_8 FILLER_10_585 ();
 sg13g2_decap_8 FILLER_10_592 ();
 sg13g2_decap_8 FILLER_10_599 ();
 sg13g2_decap_8 FILLER_10_606 ();
 sg13g2_decap_8 FILLER_10_613 ();
 sg13g2_decap_8 FILLER_10_620 ();
 sg13g2_decap_8 FILLER_10_627 ();
 sg13g2_decap_8 FILLER_10_634 ();
 sg13g2_decap_8 FILLER_10_641 ();
 sg13g2_decap_8 FILLER_10_648 ();
 sg13g2_decap_8 FILLER_10_655 ();
 sg13g2_decap_8 FILLER_10_662 ();
 sg13g2_decap_8 FILLER_10_669 ();
 sg13g2_decap_8 FILLER_10_676 ();
 sg13g2_decap_8 FILLER_10_683 ();
 sg13g2_decap_8 FILLER_10_690 ();
 sg13g2_decap_8 FILLER_10_697 ();
 sg13g2_decap_8 FILLER_10_704 ();
 sg13g2_decap_8 FILLER_10_711 ();
 sg13g2_decap_8 FILLER_10_718 ();
 sg13g2_decap_8 FILLER_10_725 ();
 sg13g2_decap_8 FILLER_10_732 ();
 sg13g2_decap_8 FILLER_10_739 ();
 sg13g2_decap_8 FILLER_10_746 ();
 sg13g2_decap_8 FILLER_10_753 ();
 sg13g2_decap_8 FILLER_10_760 ();
 sg13g2_decap_8 FILLER_10_767 ();
 sg13g2_decap_8 FILLER_10_774 ();
 sg13g2_decap_8 FILLER_10_781 ();
 sg13g2_decap_8 FILLER_10_788 ();
 sg13g2_decap_8 FILLER_10_795 ();
 sg13g2_decap_8 FILLER_10_802 ();
 sg13g2_decap_8 FILLER_10_809 ();
 sg13g2_decap_8 FILLER_10_816 ();
 sg13g2_decap_8 FILLER_10_823 ();
 sg13g2_decap_8 FILLER_10_830 ();
 sg13g2_decap_8 FILLER_10_837 ();
 sg13g2_decap_8 FILLER_10_844 ();
 sg13g2_decap_8 FILLER_10_851 ();
 sg13g2_decap_8 FILLER_10_858 ();
 sg13g2_decap_8 FILLER_10_865 ();
 sg13g2_decap_8 FILLER_10_872 ();
 sg13g2_decap_8 FILLER_10_879 ();
 sg13g2_decap_8 FILLER_10_886 ();
 sg13g2_decap_8 FILLER_10_893 ();
 sg13g2_decap_8 FILLER_10_900 ();
 sg13g2_decap_8 FILLER_10_907 ();
 sg13g2_decap_8 FILLER_10_914 ();
 sg13g2_decap_8 FILLER_10_921 ();
 sg13g2_decap_8 FILLER_10_928 ();
 sg13g2_decap_8 FILLER_10_935 ();
 sg13g2_decap_8 FILLER_10_942 ();
 sg13g2_decap_8 FILLER_10_949 ();
 sg13g2_decap_8 FILLER_10_956 ();
 sg13g2_decap_8 FILLER_10_963 ();
 sg13g2_decap_8 FILLER_10_970 ();
 sg13g2_decap_8 FILLER_10_977 ();
 sg13g2_decap_8 FILLER_10_984 ();
 sg13g2_decap_8 FILLER_10_991 ();
 sg13g2_decap_8 FILLER_10_998 ();
 sg13g2_decap_8 FILLER_10_1005 ();
 sg13g2_decap_8 FILLER_10_1012 ();
 sg13g2_decap_8 FILLER_10_1019 ();
 sg13g2_fill_2 FILLER_10_1026 ();
 sg13g2_fill_1 FILLER_10_1028 ();
 sg13g2_decap_8 FILLER_11_4 ();
 sg13g2_decap_8 FILLER_11_11 ();
 sg13g2_decap_8 FILLER_11_18 ();
 sg13g2_decap_8 FILLER_11_25 ();
 sg13g2_decap_8 FILLER_11_32 ();
 sg13g2_decap_8 FILLER_11_39 ();
 sg13g2_decap_8 FILLER_11_46 ();
 sg13g2_decap_8 FILLER_11_53 ();
 sg13g2_decap_8 FILLER_11_60 ();
 sg13g2_decap_8 FILLER_11_67 ();
 sg13g2_decap_8 FILLER_11_74 ();
 sg13g2_decap_8 FILLER_11_81 ();
 sg13g2_decap_8 FILLER_11_88 ();
 sg13g2_decap_8 FILLER_11_95 ();
 sg13g2_decap_8 FILLER_11_102 ();
 sg13g2_decap_8 FILLER_11_109 ();
 sg13g2_decap_8 FILLER_11_116 ();
 sg13g2_decap_8 FILLER_11_123 ();
 sg13g2_decap_8 FILLER_11_130 ();
 sg13g2_decap_8 FILLER_11_137 ();
 sg13g2_decap_8 FILLER_11_144 ();
 sg13g2_decap_8 FILLER_11_151 ();
 sg13g2_decap_8 FILLER_11_158 ();
 sg13g2_decap_8 FILLER_11_165 ();
 sg13g2_decap_8 FILLER_11_172 ();
 sg13g2_decap_8 FILLER_11_179 ();
 sg13g2_decap_8 FILLER_11_186 ();
 sg13g2_decap_8 FILLER_11_193 ();
 sg13g2_decap_8 FILLER_11_200 ();
 sg13g2_decap_8 FILLER_11_207 ();
 sg13g2_decap_8 FILLER_11_214 ();
 sg13g2_decap_8 FILLER_11_221 ();
 sg13g2_decap_8 FILLER_11_228 ();
 sg13g2_decap_8 FILLER_11_235 ();
 sg13g2_decap_8 FILLER_11_242 ();
 sg13g2_decap_8 FILLER_11_249 ();
 sg13g2_decap_8 FILLER_11_256 ();
 sg13g2_decap_8 FILLER_11_263 ();
 sg13g2_decap_8 FILLER_11_270 ();
 sg13g2_decap_8 FILLER_11_277 ();
 sg13g2_decap_8 FILLER_11_284 ();
 sg13g2_decap_8 FILLER_11_291 ();
 sg13g2_decap_8 FILLER_11_298 ();
 sg13g2_decap_8 FILLER_11_305 ();
 sg13g2_decap_8 FILLER_11_312 ();
 sg13g2_decap_8 FILLER_11_319 ();
 sg13g2_decap_8 FILLER_11_326 ();
 sg13g2_decap_8 FILLER_11_333 ();
 sg13g2_decap_8 FILLER_11_340 ();
 sg13g2_decap_8 FILLER_11_347 ();
 sg13g2_decap_8 FILLER_11_354 ();
 sg13g2_decap_8 FILLER_11_361 ();
 sg13g2_decap_8 FILLER_11_368 ();
 sg13g2_decap_8 FILLER_11_375 ();
 sg13g2_decap_8 FILLER_11_382 ();
 sg13g2_decap_8 FILLER_11_389 ();
 sg13g2_decap_8 FILLER_11_396 ();
 sg13g2_decap_8 FILLER_11_403 ();
 sg13g2_decap_8 FILLER_11_410 ();
 sg13g2_decap_8 FILLER_11_417 ();
 sg13g2_decap_8 FILLER_11_424 ();
 sg13g2_decap_8 FILLER_11_431 ();
 sg13g2_decap_8 FILLER_11_438 ();
 sg13g2_decap_8 FILLER_11_445 ();
 sg13g2_decap_8 FILLER_11_452 ();
 sg13g2_decap_8 FILLER_11_459 ();
 sg13g2_decap_8 FILLER_11_466 ();
 sg13g2_decap_8 FILLER_11_473 ();
 sg13g2_decap_8 FILLER_11_480 ();
 sg13g2_decap_8 FILLER_11_487 ();
 sg13g2_decap_8 FILLER_11_494 ();
 sg13g2_decap_8 FILLER_11_501 ();
 sg13g2_decap_8 FILLER_11_508 ();
 sg13g2_decap_8 FILLER_11_515 ();
 sg13g2_decap_8 FILLER_11_522 ();
 sg13g2_decap_8 FILLER_11_529 ();
 sg13g2_decap_8 FILLER_11_536 ();
 sg13g2_decap_8 FILLER_11_543 ();
 sg13g2_decap_8 FILLER_11_550 ();
 sg13g2_decap_8 FILLER_11_557 ();
 sg13g2_decap_8 FILLER_11_564 ();
 sg13g2_decap_8 FILLER_11_571 ();
 sg13g2_decap_8 FILLER_11_578 ();
 sg13g2_decap_8 FILLER_11_585 ();
 sg13g2_decap_8 FILLER_11_592 ();
 sg13g2_decap_8 FILLER_11_599 ();
 sg13g2_decap_8 FILLER_11_606 ();
 sg13g2_decap_8 FILLER_11_613 ();
 sg13g2_decap_8 FILLER_11_620 ();
 sg13g2_decap_8 FILLER_11_627 ();
 sg13g2_decap_8 FILLER_11_634 ();
 sg13g2_decap_8 FILLER_11_641 ();
 sg13g2_decap_8 FILLER_11_648 ();
 sg13g2_decap_8 FILLER_11_655 ();
 sg13g2_decap_8 FILLER_11_662 ();
 sg13g2_decap_8 FILLER_11_669 ();
 sg13g2_decap_8 FILLER_11_676 ();
 sg13g2_decap_8 FILLER_11_683 ();
 sg13g2_decap_8 FILLER_11_690 ();
 sg13g2_decap_8 FILLER_11_697 ();
 sg13g2_decap_8 FILLER_11_704 ();
 sg13g2_decap_8 FILLER_11_711 ();
 sg13g2_decap_8 FILLER_11_718 ();
 sg13g2_decap_8 FILLER_11_725 ();
 sg13g2_decap_8 FILLER_11_732 ();
 sg13g2_decap_8 FILLER_11_739 ();
 sg13g2_decap_8 FILLER_11_746 ();
 sg13g2_decap_8 FILLER_11_753 ();
 sg13g2_decap_8 FILLER_11_760 ();
 sg13g2_decap_8 FILLER_11_767 ();
 sg13g2_decap_8 FILLER_11_774 ();
 sg13g2_decap_8 FILLER_11_781 ();
 sg13g2_decap_8 FILLER_11_788 ();
 sg13g2_decap_8 FILLER_11_795 ();
 sg13g2_decap_8 FILLER_11_802 ();
 sg13g2_decap_8 FILLER_11_809 ();
 sg13g2_decap_8 FILLER_11_816 ();
 sg13g2_decap_8 FILLER_11_823 ();
 sg13g2_decap_8 FILLER_11_830 ();
 sg13g2_decap_8 FILLER_11_837 ();
 sg13g2_decap_8 FILLER_11_844 ();
 sg13g2_decap_8 FILLER_11_851 ();
 sg13g2_decap_8 FILLER_11_858 ();
 sg13g2_decap_8 FILLER_11_865 ();
 sg13g2_decap_8 FILLER_11_872 ();
 sg13g2_decap_8 FILLER_11_879 ();
 sg13g2_decap_8 FILLER_11_886 ();
 sg13g2_decap_8 FILLER_11_893 ();
 sg13g2_decap_8 FILLER_11_900 ();
 sg13g2_decap_8 FILLER_11_907 ();
 sg13g2_decap_8 FILLER_11_914 ();
 sg13g2_decap_8 FILLER_11_921 ();
 sg13g2_decap_8 FILLER_11_928 ();
 sg13g2_decap_8 FILLER_11_935 ();
 sg13g2_decap_8 FILLER_11_942 ();
 sg13g2_decap_8 FILLER_11_949 ();
 sg13g2_decap_8 FILLER_11_956 ();
 sg13g2_decap_8 FILLER_11_963 ();
 sg13g2_decap_8 FILLER_11_970 ();
 sg13g2_decap_8 FILLER_11_977 ();
 sg13g2_decap_8 FILLER_11_984 ();
 sg13g2_decap_8 FILLER_11_991 ();
 sg13g2_decap_8 FILLER_11_998 ();
 sg13g2_decap_8 FILLER_11_1005 ();
 sg13g2_decap_8 FILLER_11_1012 ();
 sg13g2_decap_8 FILLER_11_1019 ();
 sg13g2_fill_2 FILLER_11_1026 ();
 sg13g2_fill_1 FILLER_11_1028 ();
 sg13g2_decap_8 FILLER_12_4 ();
 sg13g2_decap_8 FILLER_12_11 ();
 sg13g2_decap_8 FILLER_12_18 ();
 sg13g2_decap_8 FILLER_12_25 ();
 sg13g2_decap_8 FILLER_12_32 ();
 sg13g2_decap_8 FILLER_12_39 ();
 sg13g2_decap_8 FILLER_12_46 ();
 sg13g2_decap_8 FILLER_12_53 ();
 sg13g2_decap_8 FILLER_12_60 ();
 sg13g2_decap_8 FILLER_12_67 ();
 sg13g2_decap_8 FILLER_12_74 ();
 sg13g2_decap_8 FILLER_12_81 ();
 sg13g2_decap_8 FILLER_12_88 ();
 sg13g2_decap_8 FILLER_12_95 ();
 sg13g2_decap_8 FILLER_12_102 ();
 sg13g2_decap_8 FILLER_12_109 ();
 sg13g2_decap_8 FILLER_12_116 ();
 sg13g2_decap_8 FILLER_12_123 ();
 sg13g2_decap_8 FILLER_12_130 ();
 sg13g2_decap_8 FILLER_12_137 ();
 sg13g2_decap_8 FILLER_12_144 ();
 sg13g2_decap_8 FILLER_12_151 ();
 sg13g2_decap_8 FILLER_12_158 ();
 sg13g2_decap_8 FILLER_12_165 ();
 sg13g2_decap_8 FILLER_12_172 ();
 sg13g2_decap_8 FILLER_12_179 ();
 sg13g2_decap_8 FILLER_12_186 ();
 sg13g2_decap_8 FILLER_12_193 ();
 sg13g2_decap_8 FILLER_12_200 ();
 sg13g2_decap_8 FILLER_12_207 ();
 sg13g2_decap_8 FILLER_12_214 ();
 sg13g2_decap_8 FILLER_12_221 ();
 sg13g2_decap_8 FILLER_12_228 ();
 sg13g2_decap_8 FILLER_12_235 ();
 sg13g2_decap_8 FILLER_12_242 ();
 sg13g2_decap_8 FILLER_12_249 ();
 sg13g2_decap_8 FILLER_12_256 ();
 sg13g2_decap_8 FILLER_12_263 ();
 sg13g2_decap_8 FILLER_12_270 ();
 sg13g2_decap_8 FILLER_12_277 ();
 sg13g2_decap_8 FILLER_12_284 ();
 sg13g2_decap_8 FILLER_12_291 ();
 sg13g2_decap_8 FILLER_12_298 ();
 sg13g2_decap_8 FILLER_12_305 ();
 sg13g2_decap_8 FILLER_12_312 ();
 sg13g2_decap_8 FILLER_12_319 ();
 sg13g2_decap_8 FILLER_12_326 ();
 sg13g2_decap_8 FILLER_12_333 ();
 sg13g2_decap_8 FILLER_12_340 ();
 sg13g2_decap_8 FILLER_12_347 ();
 sg13g2_decap_8 FILLER_12_354 ();
 sg13g2_decap_8 FILLER_12_361 ();
 sg13g2_decap_8 FILLER_12_368 ();
 sg13g2_decap_8 FILLER_12_375 ();
 sg13g2_decap_8 FILLER_12_382 ();
 sg13g2_decap_8 FILLER_12_389 ();
 sg13g2_decap_8 FILLER_12_396 ();
 sg13g2_decap_8 FILLER_12_403 ();
 sg13g2_decap_8 FILLER_12_410 ();
 sg13g2_decap_8 FILLER_12_417 ();
 sg13g2_decap_8 FILLER_12_424 ();
 sg13g2_decap_8 FILLER_12_431 ();
 sg13g2_decap_8 FILLER_12_438 ();
 sg13g2_decap_8 FILLER_12_445 ();
 sg13g2_decap_8 FILLER_12_452 ();
 sg13g2_decap_8 FILLER_12_459 ();
 sg13g2_decap_8 FILLER_12_466 ();
 sg13g2_decap_8 FILLER_12_473 ();
 sg13g2_decap_8 FILLER_12_480 ();
 sg13g2_decap_8 FILLER_12_487 ();
 sg13g2_decap_8 FILLER_12_494 ();
 sg13g2_decap_8 FILLER_12_501 ();
 sg13g2_decap_8 FILLER_12_508 ();
 sg13g2_decap_8 FILLER_12_515 ();
 sg13g2_decap_8 FILLER_12_522 ();
 sg13g2_decap_8 FILLER_12_529 ();
 sg13g2_decap_8 FILLER_12_536 ();
 sg13g2_decap_8 FILLER_12_543 ();
 sg13g2_decap_8 FILLER_12_550 ();
 sg13g2_decap_8 FILLER_12_557 ();
 sg13g2_decap_8 FILLER_12_564 ();
 sg13g2_decap_8 FILLER_12_571 ();
 sg13g2_decap_8 FILLER_12_578 ();
 sg13g2_decap_8 FILLER_12_585 ();
 sg13g2_decap_8 FILLER_12_592 ();
 sg13g2_decap_8 FILLER_12_599 ();
 sg13g2_decap_8 FILLER_12_606 ();
 sg13g2_decap_8 FILLER_12_613 ();
 sg13g2_decap_8 FILLER_12_620 ();
 sg13g2_decap_8 FILLER_12_627 ();
 sg13g2_decap_8 FILLER_12_634 ();
 sg13g2_decap_8 FILLER_12_641 ();
 sg13g2_decap_8 FILLER_12_648 ();
 sg13g2_decap_8 FILLER_12_655 ();
 sg13g2_decap_8 FILLER_12_662 ();
 sg13g2_decap_8 FILLER_12_669 ();
 sg13g2_decap_8 FILLER_12_676 ();
 sg13g2_decap_8 FILLER_12_683 ();
 sg13g2_decap_8 FILLER_12_690 ();
 sg13g2_decap_8 FILLER_12_697 ();
 sg13g2_decap_8 FILLER_12_704 ();
 sg13g2_decap_8 FILLER_12_711 ();
 sg13g2_decap_8 FILLER_12_718 ();
 sg13g2_decap_8 FILLER_12_725 ();
 sg13g2_decap_8 FILLER_12_732 ();
 sg13g2_decap_8 FILLER_12_739 ();
 sg13g2_decap_8 FILLER_12_746 ();
 sg13g2_decap_8 FILLER_12_753 ();
 sg13g2_decap_8 FILLER_12_760 ();
 sg13g2_decap_8 FILLER_12_767 ();
 sg13g2_decap_8 FILLER_12_774 ();
 sg13g2_decap_8 FILLER_12_781 ();
 sg13g2_decap_8 FILLER_12_788 ();
 sg13g2_decap_8 FILLER_12_795 ();
 sg13g2_decap_8 FILLER_12_802 ();
 sg13g2_decap_8 FILLER_12_809 ();
 sg13g2_decap_8 FILLER_12_816 ();
 sg13g2_decap_8 FILLER_12_823 ();
 sg13g2_decap_8 FILLER_12_830 ();
 sg13g2_decap_8 FILLER_12_837 ();
 sg13g2_decap_8 FILLER_12_844 ();
 sg13g2_decap_8 FILLER_12_851 ();
 sg13g2_decap_8 FILLER_12_858 ();
 sg13g2_decap_8 FILLER_12_865 ();
 sg13g2_decap_8 FILLER_12_872 ();
 sg13g2_decap_8 FILLER_12_879 ();
 sg13g2_decap_8 FILLER_12_886 ();
 sg13g2_decap_8 FILLER_12_893 ();
 sg13g2_decap_8 FILLER_12_900 ();
 sg13g2_decap_8 FILLER_12_907 ();
 sg13g2_decap_8 FILLER_12_914 ();
 sg13g2_decap_8 FILLER_12_921 ();
 sg13g2_decap_8 FILLER_12_928 ();
 sg13g2_decap_8 FILLER_12_935 ();
 sg13g2_decap_8 FILLER_12_942 ();
 sg13g2_decap_8 FILLER_12_949 ();
 sg13g2_decap_8 FILLER_12_956 ();
 sg13g2_decap_8 FILLER_12_963 ();
 sg13g2_decap_8 FILLER_12_970 ();
 sg13g2_decap_8 FILLER_12_977 ();
 sg13g2_decap_8 FILLER_12_984 ();
 sg13g2_decap_8 FILLER_12_991 ();
 sg13g2_decap_8 FILLER_12_998 ();
 sg13g2_decap_8 FILLER_12_1005 ();
 sg13g2_decap_8 FILLER_12_1012 ();
 sg13g2_decap_8 FILLER_12_1019 ();
 sg13g2_fill_2 FILLER_12_1026 ();
 sg13g2_fill_1 FILLER_12_1028 ();
 sg13g2_decap_8 FILLER_13_4 ();
 sg13g2_decap_8 FILLER_13_11 ();
 sg13g2_decap_8 FILLER_13_18 ();
 sg13g2_decap_8 FILLER_13_25 ();
 sg13g2_decap_8 FILLER_13_32 ();
 sg13g2_decap_8 FILLER_13_39 ();
 sg13g2_decap_8 FILLER_13_46 ();
 sg13g2_decap_8 FILLER_13_53 ();
 sg13g2_decap_8 FILLER_13_60 ();
 sg13g2_decap_8 FILLER_13_67 ();
 sg13g2_decap_8 FILLER_13_74 ();
 sg13g2_decap_8 FILLER_13_81 ();
 sg13g2_decap_8 FILLER_13_88 ();
 sg13g2_decap_8 FILLER_13_95 ();
 sg13g2_decap_8 FILLER_13_102 ();
 sg13g2_decap_8 FILLER_13_109 ();
 sg13g2_decap_8 FILLER_13_116 ();
 sg13g2_decap_8 FILLER_13_123 ();
 sg13g2_decap_8 FILLER_13_130 ();
 sg13g2_decap_8 FILLER_13_137 ();
 sg13g2_decap_8 FILLER_13_144 ();
 sg13g2_decap_8 FILLER_13_151 ();
 sg13g2_decap_8 FILLER_13_158 ();
 sg13g2_decap_8 FILLER_13_165 ();
 sg13g2_decap_8 FILLER_13_172 ();
 sg13g2_decap_8 FILLER_13_179 ();
 sg13g2_decap_8 FILLER_13_186 ();
 sg13g2_decap_8 FILLER_13_193 ();
 sg13g2_decap_8 FILLER_13_200 ();
 sg13g2_decap_8 FILLER_13_207 ();
 sg13g2_decap_8 FILLER_13_214 ();
 sg13g2_decap_8 FILLER_13_221 ();
 sg13g2_decap_8 FILLER_13_228 ();
 sg13g2_decap_8 FILLER_13_235 ();
 sg13g2_decap_8 FILLER_13_242 ();
 sg13g2_decap_8 FILLER_13_249 ();
 sg13g2_decap_8 FILLER_13_256 ();
 sg13g2_decap_8 FILLER_13_263 ();
 sg13g2_decap_8 FILLER_13_270 ();
 sg13g2_decap_8 FILLER_13_277 ();
 sg13g2_decap_8 FILLER_13_284 ();
 sg13g2_decap_8 FILLER_13_291 ();
 sg13g2_decap_8 FILLER_13_298 ();
 sg13g2_decap_8 FILLER_13_305 ();
 sg13g2_decap_8 FILLER_13_312 ();
 sg13g2_decap_8 FILLER_13_319 ();
 sg13g2_decap_8 FILLER_13_326 ();
 sg13g2_decap_8 FILLER_13_333 ();
 sg13g2_decap_8 FILLER_13_340 ();
 sg13g2_decap_8 FILLER_13_347 ();
 sg13g2_decap_8 FILLER_13_354 ();
 sg13g2_decap_8 FILLER_13_361 ();
 sg13g2_decap_8 FILLER_13_368 ();
 sg13g2_decap_8 FILLER_13_375 ();
 sg13g2_decap_8 FILLER_13_382 ();
 sg13g2_decap_8 FILLER_13_389 ();
 sg13g2_decap_8 FILLER_13_396 ();
 sg13g2_decap_8 FILLER_13_403 ();
 sg13g2_decap_8 FILLER_13_410 ();
 sg13g2_decap_8 FILLER_13_417 ();
 sg13g2_decap_8 FILLER_13_424 ();
 sg13g2_decap_8 FILLER_13_431 ();
 sg13g2_decap_8 FILLER_13_438 ();
 sg13g2_decap_8 FILLER_13_445 ();
 sg13g2_decap_8 FILLER_13_452 ();
 sg13g2_decap_8 FILLER_13_459 ();
 sg13g2_decap_8 FILLER_13_466 ();
 sg13g2_decap_8 FILLER_13_473 ();
 sg13g2_decap_8 FILLER_13_480 ();
 sg13g2_decap_8 FILLER_13_487 ();
 sg13g2_decap_8 FILLER_13_494 ();
 sg13g2_decap_8 FILLER_13_501 ();
 sg13g2_decap_8 FILLER_13_508 ();
 sg13g2_decap_8 FILLER_13_515 ();
 sg13g2_decap_8 FILLER_13_522 ();
 sg13g2_decap_8 FILLER_13_529 ();
 sg13g2_decap_8 FILLER_13_536 ();
 sg13g2_decap_8 FILLER_13_543 ();
 sg13g2_decap_8 FILLER_13_550 ();
 sg13g2_decap_8 FILLER_13_557 ();
 sg13g2_decap_8 FILLER_13_564 ();
 sg13g2_decap_8 FILLER_13_571 ();
 sg13g2_decap_8 FILLER_13_578 ();
 sg13g2_decap_8 FILLER_13_585 ();
 sg13g2_decap_8 FILLER_13_592 ();
 sg13g2_decap_8 FILLER_13_599 ();
 sg13g2_decap_8 FILLER_13_606 ();
 sg13g2_decap_8 FILLER_13_613 ();
 sg13g2_decap_8 FILLER_13_620 ();
 sg13g2_decap_8 FILLER_13_627 ();
 sg13g2_decap_8 FILLER_13_634 ();
 sg13g2_decap_8 FILLER_13_641 ();
 sg13g2_decap_8 FILLER_13_648 ();
 sg13g2_decap_8 FILLER_13_655 ();
 sg13g2_decap_8 FILLER_13_662 ();
 sg13g2_decap_8 FILLER_13_669 ();
 sg13g2_decap_8 FILLER_13_676 ();
 sg13g2_decap_8 FILLER_13_683 ();
 sg13g2_decap_8 FILLER_13_690 ();
 sg13g2_decap_8 FILLER_13_697 ();
 sg13g2_decap_8 FILLER_13_704 ();
 sg13g2_decap_8 FILLER_13_711 ();
 sg13g2_decap_8 FILLER_13_718 ();
 sg13g2_decap_8 FILLER_13_725 ();
 sg13g2_decap_8 FILLER_13_732 ();
 sg13g2_decap_8 FILLER_13_739 ();
 sg13g2_decap_8 FILLER_13_746 ();
 sg13g2_decap_8 FILLER_13_753 ();
 sg13g2_decap_8 FILLER_13_760 ();
 sg13g2_decap_8 FILLER_13_767 ();
 sg13g2_decap_8 FILLER_13_774 ();
 sg13g2_decap_8 FILLER_13_781 ();
 sg13g2_decap_8 FILLER_13_788 ();
 sg13g2_decap_8 FILLER_13_795 ();
 sg13g2_decap_8 FILLER_13_802 ();
 sg13g2_decap_8 FILLER_13_809 ();
 sg13g2_decap_8 FILLER_13_816 ();
 sg13g2_decap_8 FILLER_13_823 ();
 sg13g2_decap_8 FILLER_13_830 ();
 sg13g2_decap_8 FILLER_13_837 ();
 sg13g2_decap_8 FILLER_13_844 ();
 sg13g2_decap_8 FILLER_13_851 ();
 sg13g2_decap_8 FILLER_13_858 ();
 sg13g2_decap_8 FILLER_13_865 ();
 sg13g2_decap_8 FILLER_13_872 ();
 sg13g2_decap_8 FILLER_13_879 ();
 sg13g2_decap_8 FILLER_13_886 ();
 sg13g2_decap_8 FILLER_13_893 ();
 sg13g2_decap_8 FILLER_13_900 ();
 sg13g2_decap_8 FILLER_13_907 ();
 sg13g2_decap_8 FILLER_13_914 ();
 sg13g2_decap_8 FILLER_13_921 ();
 sg13g2_decap_8 FILLER_13_928 ();
 sg13g2_decap_8 FILLER_13_935 ();
 sg13g2_decap_8 FILLER_13_942 ();
 sg13g2_decap_8 FILLER_13_949 ();
 sg13g2_decap_8 FILLER_13_956 ();
 sg13g2_decap_8 FILLER_13_963 ();
 sg13g2_decap_8 FILLER_13_970 ();
 sg13g2_decap_8 FILLER_13_977 ();
 sg13g2_decap_8 FILLER_13_984 ();
 sg13g2_decap_8 FILLER_13_991 ();
 sg13g2_decap_8 FILLER_13_998 ();
 sg13g2_decap_8 FILLER_13_1005 ();
 sg13g2_decap_8 FILLER_13_1012 ();
 sg13g2_decap_8 FILLER_13_1019 ();
 sg13g2_fill_2 FILLER_13_1026 ();
 sg13g2_fill_1 FILLER_13_1028 ();
 sg13g2_decap_8 FILLER_14_4 ();
 sg13g2_decap_8 FILLER_14_11 ();
 sg13g2_decap_8 FILLER_14_18 ();
 sg13g2_decap_8 FILLER_14_25 ();
 sg13g2_decap_8 FILLER_14_32 ();
 sg13g2_decap_8 FILLER_14_39 ();
 sg13g2_decap_8 FILLER_14_46 ();
 sg13g2_decap_8 FILLER_14_53 ();
 sg13g2_decap_8 FILLER_14_60 ();
 sg13g2_decap_8 FILLER_14_67 ();
 sg13g2_decap_8 FILLER_14_74 ();
 sg13g2_decap_8 FILLER_14_81 ();
 sg13g2_decap_8 FILLER_14_88 ();
 sg13g2_decap_8 FILLER_14_95 ();
 sg13g2_decap_8 FILLER_14_102 ();
 sg13g2_decap_8 FILLER_14_109 ();
 sg13g2_decap_8 FILLER_14_116 ();
 sg13g2_decap_8 FILLER_14_123 ();
 sg13g2_decap_8 FILLER_14_130 ();
 sg13g2_decap_8 FILLER_14_137 ();
 sg13g2_decap_8 FILLER_14_144 ();
 sg13g2_decap_8 FILLER_14_151 ();
 sg13g2_decap_8 FILLER_14_158 ();
 sg13g2_decap_8 FILLER_14_165 ();
 sg13g2_decap_8 FILLER_14_172 ();
 sg13g2_decap_8 FILLER_14_179 ();
 sg13g2_decap_8 FILLER_14_186 ();
 sg13g2_decap_8 FILLER_14_193 ();
 sg13g2_decap_8 FILLER_14_200 ();
 sg13g2_decap_8 FILLER_14_207 ();
 sg13g2_decap_8 FILLER_14_214 ();
 sg13g2_decap_8 FILLER_14_221 ();
 sg13g2_decap_8 FILLER_14_255 ();
 sg13g2_decap_8 FILLER_14_262 ();
 sg13g2_decap_8 FILLER_14_269 ();
 sg13g2_decap_8 FILLER_14_276 ();
 sg13g2_decap_8 FILLER_14_283 ();
 sg13g2_decap_8 FILLER_14_290 ();
 sg13g2_decap_8 FILLER_14_297 ();
 sg13g2_decap_8 FILLER_14_304 ();
 sg13g2_decap_8 FILLER_14_311 ();
 sg13g2_decap_8 FILLER_14_318 ();
 sg13g2_decap_8 FILLER_14_325 ();
 sg13g2_decap_8 FILLER_14_332 ();
 sg13g2_decap_8 FILLER_14_339 ();
 sg13g2_decap_8 FILLER_14_346 ();
 sg13g2_decap_8 FILLER_14_353 ();
 sg13g2_decap_8 FILLER_14_360 ();
 sg13g2_decap_8 FILLER_14_367 ();
 sg13g2_decap_8 FILLER_14_374 ();
 sg13g2_decap_8 FILLER_14_381 ();
 sg13g2_decap_8 FILLER_14_388 ();
 sg13g2_decap_8 FILLER_14_395 ();
 sg13g2_decap_8 FILLER_14_402 ();
 sg13g2_decap_8 FILLER_14_409 ();
 sg13g2_decap_8 FILLER_14_416 ();
 sg13g2_decap_8 FILLER_14_423 ();
 sg13g2_decap_8 FILLER_14_430 ();
 sg13g2_decap_8 FILLER_14_437 ();
 sg13g2_decap_8 FILLER_14_444 ();
 sg13g2_decap_8 FILLER_14_451 ();
 sg13g2_decap_8 FILLER_14_458 ();
 sg13g2_decap_8 FILLER_14_465 ();
 sg13g2_decap_8 FILLER_14_472 ();
 sg13g2_decap_8 FILLER_14_479 ();
 sg13g2_decap_8 FILLER_14_486 ();
 sg13g2_decap_8 FILLER_14_493 ();
 sg13g2_decap_8 FILLER_14_500 ();
 sg13g2_decap_8 FILLER_14_507 ();
 sg13g2_decap_8 FILLER_14_514 ();
 sg13g2_decap_8 FILLER_14_521 ();
 sg13g2_decap_8 FILLER_14_528 ();
 sg13g2_decap_8 FILLER_14_535 ();
 sg13g2_decap_8 FILLER_14_542 ();
 sg13g2_decap_8 FILLER_14_549 ();
 sg13g2_decap_8 FILLER_14_556 ();
 sg13g2_decap_8 FILLER_14_563 ();
 sg13g2_decap_8 FILLER_14_570 ();
 sg13g2_decap_8 FILLER_14_577 ();
 sg13g2_decap_8 FILLER_14_584 ();
 sg13g2_decap_8 FILLER_14_591 ();
 sg13g2_decap_8 FILLER_14_598 ();
 sg13g2_decap_8 FILLER_14_605 ();
 sg13g2_decap_8 FILLER_14_612 ();
 sg13g2_decap_8 FILLER_14_619 ();
 sg13g2_decap_8 FILLER_14_626 ();
 sg13g2_decap_8 FILLER_14_633 ();
 sg13g2_decap_8 FILLER_14_640 ();
 sg13g2_decap_8 FILLER_14_647 ();
 sg13g2_decap_8 FILLER_14_654 ();
 sg13g2_decap_8 FILLER_14_661 ();
 sg13g2_decap_8 FILLER_14_668 ();
 sg13g2_decap_8 FILLER_14_675 ();
 sg13g2_decap_8 FILLER_14_682 ();
 sg13g2_decap_8 FILLER_14_689 ();
 sg13g2_decap_8 FILLER_14_696 ();
 sg13g2_decap_8 FILLER_14_703 ();
 sg13g2_decap_8 FILLER_14_710 ();
 sg13g2_decap_8 FILLER_14_717 ();
 sg13g2_decap_8 FILLER_14_724 ();
 sg13g2_decap_8 FILLER_14_731 ();
 sg13g2_decap_8 FILLER_14_738 ();
 sg13g2_decap_8 FILLER_14_745 ();
 sg13g2_decap_8 FILLER_14_752 ();
 sg13g2_decap_8 FILLER_14_759 ();
 sg13g2_decap_8 FILLER_14_766 ();
 sg13g2_decap_8 FILLER_14_773 ();
 sg13g2_decap_8 FILLER_14_780 ();
 sg13g2_decap_8 FILLER_14_787 ();
 sg13g2_decap_8 FILLER_14_794 ();
 sg13g2_decap_8 FILLER_14_801 ();
 sg13g2_decap_8 FILLER_14_808 ();
 sg13g2_decap_8 FILLER_14_815 ();
 sg13g2_decap_8 FILLER_14_822 ();
 sg13g2_decap_8 FILLER_14_829 ();
 sg13g2_decap_8 FILLER_14_836 ();
 sg13g2_decap_8 FILLER_14_843 ();
 sg13g2_decap_8 FILLER_14_850 ();
 sg13g2_decap_8 FILLER_14_857 ();
 sg13g2_decap_8 FILLER_14_864 ();
 sg13g2_decap_8 FILLER_14_871 ();
 sg13g2_decap_8 FILLER_14_878 ();
 sg13g2_decap_8 FILLER_14_885 ();
 sg13g2_decap_8 FILLER_14_892 ();
 sg13g2_decap_8 FILLER_14_899 ();
 sg13g2_decap_8 FILLER_14_906 ();
 sg13g2_decap_8 FILLER_14_913 ();
 sg13g2_decap_8 FILLER_14_920 ();
 sg13g2_decap_8 FILLER_14_927 ();
 sg13g2_decap_8 FILLER_14_934 ();
 sg13g2_decap_8 FILLER_14_941 ();
 sg13g2_decap_8 FILLER_14_948 ();
 sg13g2_decap_8 FILLER_14_955 ();
 sg13g2_decap_8 FILLER_14_962 ();
 sg13g2_decap_8 FILLER_14_969 ();
 sg13g2_decap_8 FILLER_14_976 ();
 sg13g2_decap_8 FILLER_14_983 ();
 sg13g2_decap_8 FILLER_14_990 ();
 sg13g2_decap_8 FILLER_14_997 ();
 sg13g2_decap_8 FILLER_14_1004 ();
 sg13g2_decap_8 FILLER_14_1011 ();
 sg13g2_decap_8 FILLER_14_1018 ();
 sg13g2_decap_4 FILLER_14_1025 ();
 sg13g2_decap_8 FILLER_15_4 ();
 sg13g2_decap_8 FILLER_15_11 ();
 sg13g2_decap_8 FILLER_15_18 ();
 sg13g2_decap_8 FILLER_15_25 ();
 sg13g2_decap_8 FILLER_15_32 ();
 sg13g2_decap_8 FILLER_15_39 ();
 sg13g2_decap_8 FILLER_15_46 ();
 sg13g2_decap_8 FILLER_15_53 ();
 sg13g2_decap_8 FILLER_15_60 ();
 sg13g2_decap_8 FILLER_15_67 ();
 sg13g2_decap_8 FILLER_15_74 ();
 sg13g2_decap_8 FILLER_15_81 ();
 sg13g2_decap_8 FILLER_15_88 ();
 sg13g2_decap_8 FILLER_15_95 ();
 sg13g2_decap_8 FILLER_15_102 ();
 sg13g2_decap_8 FILLER_15_109 ();
 sg13g2_decap_8 FILLER_15_116 ();
 sg13g2_decap_8 FILLER_15_123 ();
 sg13g2_decap_8 FILLER_15_130 ();
 sg13g2_decap_8 FILLER_15_137 ();
 sg13g2_decap_8 FILLER_15_144 ();
 sg13g2_decap_8 FILLER_15_151 ();
 sg13g2_decap_8 FILLER_15_158 ();
 sg13g2_decap_8 FILLER_15_165 ();
 sg13g2_decap_4 FILLER_15_172 ();
 sg13g2_fill_2 FILLER_15_176 ();
 sg13g2_decap_8 FILLER_15_205 ();
 sg13g2_decap_8 FILLER_15_212 ();
 sg13g2_decap_8 FILLER_15_219 ();
 sg13g2_decap_8 FILLER_15_226 ();
 sg13g2_decap_8 FILLER_15_233 ();
 sg13g2_decap_8 FILLER_15_240 ();
 sg13g2_decap_8 FILLER_15_247 ();
 sg13g2_decap_8 FILLER_15_254 ();
 sg13g2_decap_8 FILLER_15_261 ();
 sg13g2_decap_8 FILLER_15_288 ();
 sg13g2_decap_8 FILLER_15_295 ();
 sg13g2_decap_8 FILLER_15_302 ();
 sg13g2_fill_2 FILLER_15_309 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_decap_8 FILLER_15_406 ();
 sg13g2_decap_8 FILLER_15_413 ();
 sg13g2_decap_8 FILLER_15_420 ();
 sg13g2_decap_8 FILLER_15_427 ();
 sg13g2_decap_8 FILLER_15_434 ();
 sg13g2_decap_8 FILLER_15_441 ();
 sg13g2_decap_8 FILLER_15_448 ();
 sg13g2_decap_8 FILLER_15_455 ();
 sg13g2_decap_8 FILLER_15_462 ();
 sg13g2_decap_8 FILLER_15_469 ();
 sg13g2_decap_8 FILLER_15_476 ();
 sg13g2_decap_8 FILLER_15_483 ();
 sg13g2_decap_8 FILLER_15_490 ();
 sg13g2_decap_8 FILLER_15_497 ();
 sg13g2_decap_8 FILLER_15_504 ();
 sg13g2_decap_8 FILLER_15_511 ();
 sg13g2_decap_8 FILLER_15_518 ();
 sg13g2_decap_8 FILLER_15_525 ();
 sg13g2_decap_8 FILLER_15_532 ();
 sg13g2_decap_8 FILLER_15_539 ();
 sg13g2_decap_8 FILLER_15_546 ();
 sg13g2_decap_8 FILLER_15_553 ();
 sg13g2_decap_8 FILLER_15_560 ();
 sg13g2_decap_8 FILLER_15_567 ();
 sg13g2_decap_8 FILLER_15_574 ();
 sg13g2_decap_8 FILLER_15_581 ();
 sg13g2_decap_8 FILLER_15_588 ();
 sg13g2_decap_8 FILLER_15_595 ();
 sg13g2_decap_8 FILLER_15_602 ();
 sg13g2_decap_8 FILLER_15_609 ();
 sg13g2_decap_8 FILLER_15_616 ();
 sg13g2_decap_8 FILLER_15_623 ();
 sg13g2_decap_8 FILLER_15_630 ();
 sg13g2_decap_8 FILLER_15_637 ();
 sg13g2_decap_8 FILLER_15_644 ();
 sg13g2_decap_8 FILLER_15_651 ();
 sg13g2_decap_8 FILLER_15_658 ();
 sg13g2_decap_8 FILLER_15_665 ();
 sg13g2_decap_8 FILLER_15_672 ();
 sg13g2_decap_8 FILLER_15_679 ();
 sg13g2_decap_8 FILLER_15_686 ();
 sg13g2_decap_8 FILLER_15_693 ();
 sg13g2_decap_8 FILLER_15_700 ();
 sg13g2_decap_8 FILLER_15_707 ();
 sg13g2_decap_8 FILLER_15_714 ();
 sg13g2_decap_8 FILLER_15_721 ();
 sg13g2_decap_8 FILLER_15_728 ();
 sg13g2_decap_8 FILLER_15_735 ();
 sg13g2_decap_8 FILLER_15_742 ();
 sg13g2_decap_8 FILLER_15_749 ();
 sg13g2_decap_8 FILLER_15_756 ();
 sg13g2_decap_8 FILLER_15_763 ();
 sg13g2_decap_8 FILLER_15_770 ();
 sg13g2_decap_8 FILLER_15_777 ();
 sg13g2_decap_8 FILLER_15_784 ();
 sg13g2_decap_8 FILLER_15_791 ();
 sg13g2_decap_8 FILLER_15_798 ();
 sg13g2_decap_8 FILLER_15_805 ();
 sg13g2_decap_8 FILLER_15_812 ();
 sg13g2_decap_8 FILLER_15_819 ();
 sg13g2_decap_8 FILLER_15_826 ();
 sg13g2_decap_8 FILLER_15_833 ();
 sg13g2_decap_8 FILLER_15_840 ();
 sg13g2_decap_8 FILLER_15_847 ();
 sg13g2_decap_8 FILLER_15_854 ();
 sg13g2_decap_8 FILLER_15_861 ();
 sg13g2_decap_8 FILLER_15_868 ();
 sg13g2_decap_8 FILLER_15_875 ();
 sg13g2_decap_8 FILLER_15_882 ();
 sg13g2_decap_8 FILLER_15_889 ();
 sg13g2_decap_8 FILLER_15_896 ();
 sg13g2_decap_8 FILLER_15_903 ();
 sg13g2_decap_8 FILLER_15_910 ();
 sg13g2_decap_8 FILLER_15_917 ();
 sg13g2_decap_8 FILLER_15_924 ();
 sg13g2_decap_8 FILLER_15_931 ();
 sg13g2_decap_8 FILLER_15_938 ();
 sg13g2_decap_8 FILLER_15_945 ();
 sg13g2_decap_8 FILLER_15_952 ();
 sg13g2_decap_8 FILLER_15_959 ();
 sg13g2_decap_8 FILLER_15_966 ();
 sg13g2_decap_8 FILLER_15_973 ();
 sg13g2_decap_8 FILLER_15_980 ();
 sg13g2_decap_8 FILLER_15_987 ();
 sg13g2_decap_8 FILLER_15_994 ();
 sg13g2_decap_8 FILLER_15_1001 ();
 sg13g2_decap_8 FILLER_15_1008 ();
 sg13g2_decap_8 FILLER_15_1015 ();
 sg13g2_decap_8 FILLER_15_1022 ();
 sg13g2_decap_8 FILLER_16_4 ();
 sg13g2_decap_8 FILLER_16_11 ();
 sg13g2_decap_8 FILLER_16_18 ();
 sg13g2_decap_8 FILLER_16_25 ();
 sg13g2_decap_8 FILLER_16_32 ();
 sg13g2_decap_8 FILLER_16_39 ();
 sg13g2_decap_8 FILLER_16_46 ();
 sg13g2_decap_8 FILLER_16_53 ();
 sg13g2_decap_8 FILLER_16_60 ();
 sg13g2_decap_8 FILLER_16_67 ();
 sg13g2_decap_8 FILLER_16_74 ();
 sg13g2_decap_8 FILLER_16_81 ();
 sg13g2_decap_8 FILLER_16_88 ();
 sg13g2_decap_8 FILLER_16_95 ();
 sg13g2_decap_8 FILLER_16_102 ();
 sg13g2_decap_8 FILLER_16_109 ();
 sg13g2_decap_8 FILLER_16_116 ();
 sg13g2_decap_8 FILLER_16_123 ();
 sg13g2_decap_8 FILLER_16_130 ();
 sg13g2_decap_8 FILLER_16_137 ();
 sg13g2_decap_8 FILLER_16_144 ();
 sg13g2_decap_8 FILLER_16_151 ();
 sg13g2_decap_8 FILLER_16_158 ();
 sg13g2_decap_8 FILLER_16_165 ();
 sg13g2_decap_8 FILLER_16_172 ();
 sg13g2_decap_8 FILLER_16_179 ();
 sg13g2_decap_8 FILLER_16_186 ();
 sg13g2_decap_8 FILLER_16_193 ();
 sg13g2_decap_8 FILLER_16_200 ();
 sg13g2_decap_8 FILLER_16_207 ();
 sg13g2_decap_8 FILLER_16_214 ();
 sg13g2_decap_8 FILLER_16_221 ();
 sg13g2_decap_8 FILLER_16_228 ();
 sg13g2_decap_8 FILLER_16_235 ();
 sg13g2_decap_8 FILLER_16_242 ();
 sg13g2_decap_8 FILLER_16_249 ();
 sg13g2_decap_8 FILLER_16_256 ();
 sg13g2_decap_8 FILLER_16_263 ();
 sg13g2_decap_8 FILLER_16_270 ();
 sg13g2_decap_8 FILLER_16_277 ();
 sg13g2_decap_8 FILLER_16_284 ();
 sg13g2_decap_8 FILLER_16_291 ();
 sg13g2_decap_8 FILLER_16_298 ();
 sg13g2_decap_8 FILLER_16_305 ();
 sg13g2_decap_8 FILLER_16_312 ();
 sg13g2_decap_8 FILLER_16_319 ();
 sg13g2_decap_8 FILLER_16_326 ();
 sg13g2_decap_4 FILLER_16_333 ();
 sg13g2_decap_8 FILLER_16_342 ();
 sg13g2_decap_8 FILLER_16_349 ();
 sg13g2_decap_8 FILLER_16_356 ();
 sg13g2_decap_8 FILLER_16_363 ();
 sg13g2_decap_8 FILLER_16_370 ();
 sg13g2_decap_8 FILLER_16_377 ();
 sg13g2_decap_8 FILLER_16_384 ();
 sg13g2_decap_8 FILLER_16_391 ();
 sg13g2_decap_8 FILLER_16_398 ();
 sg13g2_decap_8 FILLER_16_405 ();
 sg13g2_decap_8 FILLER_16_412 ();
 sg13g2_decap_8 FILLER_16_419 ();
 sg13g2_decap_8 FILLER_16_426 ();
 sg13g2_decap_8 FILLER_16_433 ();
 sg13g2_decap_8 FILLER_16_440 ();
 sg13g2_decap_8 FILLER_16_447 ();
 sg13g2_decap_8 FILLER_16_454 ();
 sg13g2_decap_8 FILLER_16_461 ();
 sg13g2_decap_8 FILLER_16_468 ();
 sg13g2_decap_8 FILLER_16_475 ();
 sg13g2_decap_8 FILLER_16_482 ();
 sg13g2_decap_8 FILLER_16_489 ();
 sg13g2_decap_8 FILLER_16_496 ();
 sg13g2_decap_8 FILLER_16_503 ();
 sg13g2_decap_8 FILLER_16_510 ();
 sg13g2_decap_8 FILLER_16_517 ();
 sg13g2_decap_8 FILLER_16_524 ();
 sg13g2_decap_8 FILLER_16_531 ();
 sg13g2_decap_8 FILLER_16_538 ();
 sg13g2_decap_8 FILLER_16_545 ();
 sg13g2_decap_8 FILLER_16_552 ();
 sg13g2_decap_8 FILLER_16_559 ();
 sg13g2_decap_8 FILLER_16_566 ();
 sg13g2_decap_8 FILLER_16_573 ();
 sg13g2_decap_8 FILLER_16_580 ();
 sg13g2_decap_8 FILLER_16_587 ();
 sg13g2_decap_8 FILLER_16_594 ();
 sg13g2_decap_8 FILLER_16_601 ();
 sg13g2_decap_8 FILLER_16_608 ();
 sg13g2_decap_8 FILLER_16_615 ();
 sg13g2_decap_8 FILLER_16_622 ();
 sg13g2_decap_8 FILLER_16_629 ();
 sg13g2_decap_8 FILLER_16_636 ();
 sg13g2_decap_8 FILLER_16_643 ();
 sg13g2_decap_8 FILLER_16_650 ();
 sg13g2_decap_8 FILLER_16_657 ();
 sg13g2_decap_8 FILLER_16_664 ();
 sg13g2_decap_8 FILLER_16_671 ();
 sg13g2_decap_8 FILLER_16_678 ();
 sg13g2_decap_8 FILLER_16_685 ();
 sg13g2_decap_8 FILLER_16_692 ();
 sg13g2_decap_8 FILLER_16_699 ();
 sg13g2_decap_8 FILLER_16_706 ();
 sg13g2_decap_8 FILLER_16_713 ();
 sg13g2_decap_8 FILLER_16_720 ();
 sg13g2_decap_8 FILLER_16_727 ();
 sg13g2_decap_8 FILLER_16_734 ();
 sg13g2_decap_8 FILLER_16_741 ();
 sg13g2_decap_8 FILLER_16_748 ();
 sg13g2_decap_8 FILLER_16_755 ();
 sg13g2_decap_8 FILLER_16_762 ();
 sg13g2_decap_8 FILLER_16_769 ();
 sg13g2_decap_8 FILLER_16_776 ();
 sg13g2_decap_8 FILLER_16_783 ();
 sg13g2_decap_8 FILLER_16_790 ();
 sg13g2_decap_8 FILLER_16_797 ();
 sg13g2_decap_8 FILLER_16_804 ();
 sg13g2_decap_8 FILLER_16_811 ();
 sg13g2_decap_8 FILLER_16_818 ();
 sg13g2_decap_8 FILLER_16_825 ();
 sg13g2_decap_8 FILLER_16_832 ();
 sg13g2_decap_8 FILLER_16_839 ();
 sg13g2_decap_8 FILLER_16_846 ();
 sg13g2_decap_8 FILLER_16_853 ();
 sg13g2_decap_8 FILLER_16_860 ();
 sg13g2_decap_8 FILLER_16_867 ();
 sg13g2_decap_8 FILLER_16_874 ();
 sg13g2_decap_8 FILLER_16_881 ();
 sg13g2_decap_8 FILLER_16_888 ();
 sg13g2_decap_8 FILLER_16_895 ();
 sg13g2_decap_8 FILLER_16_902 ();
 sg13g2_decap_8 FILLER_16_909 ();
 sg13g2_decap_8 FILLER_16_916 ();
 sg13g2_decap_8 FILLER_16_923 ();
 sg13g2_decap_8 FILLER_16_930 ();
 sg13g2_decap_8 FILLER_16_937 ();
 sg13g2_decap_8 FILLER_16_944 ();
 sg13g2_decap_8 FILLER_16_951 ();
 sg13g2_decap_8 FILLER_16_958 ();
 sg13g2_decap_8 FILLER_16_965 ();
 sg13g2_decap_8 FILLER_16_972 ();
 sg13g2_decap_8 FILLER_16_979 ();
 sg13g2_decap_8 FILLER_16_986 ();
 sg13g2_decap_8 FILLER_16_993 ();
 sg13g2_decap_8 FILLER_16_1000 ();
 sg13g2_decap_8 FILLER_16_1007 ();
 sg13g2_decap_8 FILLER_16_1014 ();
 sg13g2_decap_8 FILLER_16_1021 ();
 sg13g2_fill_1 FILLER_16_1028 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_decap_8 FILLER_17_406 ();
 sg13g2_decap_8 FILLER_17_413 ();
 sg13g2_decap_8 FILLER_17_420 ();
 sg13g2_decap_8 FILLER_17_427 ();
 sg13g2_decap_8 FILLER_17_434 ();
 sg13g2_decap_8 FILLER_17_441 ();
 sg13g2_decap_8 FILLER_17_448 ();
 sg13g2_decap_8 FILLER_17_455 ();
 sg13g2_decap_8 FILLER_17_462 ();
 sg13g2_decap_8 FILLER_17_469 ();
 sg13g2_decap_8 FILLER_17_476 ();
 sg13g2_decap_8 FILLER_17_483 ();
 sg13g2_decap_8 FILLER_17_490 ();
 sg13g2_decap_8 FILLER_17_497 ();
 sg13g2_decap_8 FILLER_17_504 ();
 sg13g2_decap_8 FILLER_17_511 ();
 sg13g2_decap_8 FILLER_17_518 ();
 sg13g2_decap_8 FILLER_17_525 ();
 sg13g2_decap_8 FILLER_17_532 ();
 sg13g2_decap_8 FILLER_17_539 ();
 sg13g2_decap_8 FILLER_17_546 ();
 sg13g2_decap_8 FILLER_17_553 ();
 sg13g2_decap_8 FILLER_17_560 ();
 sg13g2_decap_8 FILLER_17_567 ();
 sg13g2_decap_8 FILLER_17_574 ();
 sg13g2_decap_8 FILLER_17_581 ();
 sg13g2_decap_8 FILLER_17_588 ();
 sg13g2_decap_8 FILLER_17_595 ();
 sg13g2_decap_8 FILLER_17_602 ();
 sg13g2_decap_8 FILLER_17_609 ();
 sg13g2_decap_8 FILLER_17_616 ();
 sg13g2_decap_8 FILLER_17_623 ();
 sg13g2_decap_8 FILLER_17_630 ();
 sg13g2_decap_8 FILLER_17_637 ();
 sg13g2_decap_8 FILLER_17_644 ();
 sg13g2_decap_8 FILLER_17_651 ();
 sg13g2_decap_8 FILLER_17_658 ();
 sg13g2_decap_8 FILLER_17_665 ();
 sg13g2_decap_8 FILLER_17_672 ();
 sg13g2_decap_8 FILLER_17_679 ();
 sg13g2_decap_8 FILLER_17_686 ();
 sg13g2_decap_8 FILLER_17_693 ();
 sg13g2_decap_8 FILLER_17_700 ();
 sg13g2_decap_8 FILLER_17_707 ();
 sg13g2_decap_8 FILLER_17_714 ();
 sg13g2_decap_8 FILLER_17_721 ();
 sg13g2_decap_8 FILLER_17_728 ();
 sg13g2_decap_8 FILLER_17_735 ();
 sg13g2_decap_8 FILLER_17_742 ();
 sg13g2_decap_8 FILLER_17_749 ();
 sg13g2_decap_8 FILLER_17_756 ();
 sg13g2_decap_8 FILLER_17_763 ();
 sg13g2_decap_8 FILLER_17_770 ();
 sg13g2_decap_8 FILLER_17_777 ();
 sg13g2_decap_8 FILLER_17_784 ();
 sg13g2_decap_8 FILLER_17_791 ();
 sg13g2_decap_8 FILLER_17_798 ();
 sg13g2_decap_8 FILLER_17_805 ();
 sg13g2_decap_8 FILLER_17_812 ();
 sg13g2_decap_8 FILLER_17_819 ();
 sg13g2_decap_8 FILLER_17_826 ();
 sg13g2_decap_8 FILLER_17_833 ();
 sg13g2_decap_8 FILLER_17_840 ();
 sg13g2_decap_8 FILLER_17_847 ();
 sg13g2_decap_8 FILLER_17_854 ();
 sg13g2_decap_8 FILLER_17_861 ();
 sg13g2_decap_8 FILLER_17_868 ();
 sg13g2_decap_8 FILLER_17_875 ();
 sg13g2_decap_8 FILLER_17_882 ();
 sg13g2_decap_8 FILLER_17_889 ();
 sg13g2_decap_8 FILLER_17_896 ();
 sg13g2_decap_8 FILLER_17_903 ();
 sg13g2_decap_8 FILLER_17_910 ();
 sg13g2_decap_8 FILLER_17_917 ();
 sg13g2_decap_8 FILLER_17_924 ();
 sg13g2_decap_8 FILLER_17_931 ();
 sg13g2_decap_8 FILLER_17_938 ();
 sg13g2_decap_8 FILLER_17_945 ();
 sg13g2_decap_8 FILLER_17_952 ();
 sg13g2_decap_8 FILLER_17_959 ();
 sg13g2_decap_8 FILLER_17_966 ();
 sg13g2_decap_8 FILLER_17_973 ();
 sg13g2_decap_8 FILLER_17_980 ();
 sg13g2_decap_8 FILLER_17_987 ();
 sg13g2_decap_8 FILLER_17_994 ();
 sg13g2_decap_8 FILLER_17_1001 ();
 sg13g2_decap_8 FILLER_17_1008 ();
 sg13g2_decap_8 FILLER_17_1015 ();
 sg13g2_decap_8 FILLER_17_1022 ();
 sg13g2_decap_8 FILLER_18_4 ();
 sg13g2_decap_8 FILLER_18_11 ();
 sg13g2_decap_8 FILLER_18_18 ();
 sg13g2_decap_8 FILLER_18_25 ();
 sg13g2_decap_8 FILLER_18_32 ();
 sg13g2_decap_8 FILLER_18_39 ();
 sg13g2_decap_8 FILLER_18_46 ();
 sg13g2_decap_8 FILLER_18_53 ();
 sg13g2_decap_8 FILLER_18_60 ();
 sg13g2_decap_8 FILLER_18_67 ();
 sg13g2_decap_8 FILLER_18_74 ();
 sg13g2_decap_8 FILLER_18_81 ();
 sg13g2_decap_8 FILLER_18_88 ();
 sg13g2_decap_8 FILLER_18_95 ();
 sg13g2_decap_8 FILLER_18_102 ();
 sg13g2_decap_8 FILLER_18_109 ();
 sg13g2_decap_8 FILLER_18_116 ();
 sg13g2_decap_8 FILLER_18_123 ();
 sg13g2_decap_8 FILLER_18_130 ();
 sg13g2_decap_8 FILLER_18_137 ();
 sg13g2_decap_8 FILLER_18_144 ();
 sg13g2_decap_8 FILLER_18_151 ();
 sg13g2_decap_8 FILLER_18_158 ();
 sg13g2_decap_8 FILLER_18_165 ();
 sg13g2_decap_8 FILLER_18_172 ();
 sg13g2_decap_8 FILLER_18_179 ();
 sg13g2_decap_8 FILLER_18_186 ();
 sg13g2_decap_8 FILLER_18_193 ();
 sg13g2_decap_8 FILLER_18_200 ();
 sg13g2_decap_8 FILLER_18_207 ();
 sg13g2_decap_8 FILLER_18_214 ();
 sg13g2_decap_8 FILLER_18_221 ();
 sg13g2_fill_1 FILLER_18_228 ();
 sg13g2_decap_8 FILLER_18_256 ();
 sg13g2_decap_8 FILLER_18_263 ();
 sg13g2_decap_8 FILLER_18_270 ();
 sg13g2_decap_8 FILLER_18_277 ();
 sg13g2_decap_8 FILLER_18_284 ();
 sg13g2_decap_8 FILLER_18_291 ();
 sg13g2_decap_8 FILLER_18_298 ();
 sg13g2_decap_8 FILLER_18_305 ();
 sg13g2_decap_8 FILLER_18_312 ();
 sg13g2_decap_8 FILLER_18_319 ();
 sg13g2_decap_8 FILLER_18_326 ();
 sg13g2_decap_8 FILLER_18_333 ();
 sg13g2_decap_8 FILLER_18_340 ();
 sg13g2_decap_8 FILLER_18_347 ();
 sg13g2_decap_8 FILLER_18_354 ();
 sg13g2_decap_8 FILLER_18_361 ();
 sg13g2_decap_8 FILLER_18_368 ();
 sg13g2_decap_8 FILLER_18_375 ();
 sg13g2_decap_8 FILLER_18_382 ();
 sg13g2_decap_8 FILLER_18_389 ();
 sg13g2_decap_8 FILLER_18_396 ();
 sg13g2_decap_8 FILLER_18_403 ();
 sg13g2_decap_8 FILLER_18_410 ();
 sg13g2_decap_8 FILLER_18_417 ();
 sg13g2_decap_8 FILLER_18_424 ();
 sg13g2_decap_8 FILLER_18_431 ();
 sg13g2_decap_8 FILLER_18_438 ();
 sg13g2_decap_8 FILLER_18_445 ();
 sg13g2_decap_8 FILLER_18_452 ();
 sg13g2_decap_8 FILLER_18_459 ();
 sg13g2_decap_8 FILLER_18_466 ();
 sg13g2_decap_8 FILLER_18_473 ();
 sg13g2_decap_8 FILLER_18_480 ();
 sg13g2_decap_8 FILLER_18_487 ();
 sg13g2_decap_8 FILLER_18_494 ();
 sg13g2_decap_8 FILLER_18_501 ();
 sg13g2_decap_8 FILLER_18_508 ();
 sg13g2_decap_8 FILLER_18_515 ();
 sg13g2_decap_8 FILLER_18_522 ();
 sg13g2_decap_8 FILLER_18_529 ();
 sg13g2_decap_8 FILLER_18_536 ();
 sg13g2_decap_8 FILLER_18_543 ();
 sg13g2_decap_8 FILLER_18_550 ();
 sg13g2_decap_8 FILLER_18_557 ();
 sg13g2_decap_8 FILLER_18_564 ();
 sg13g2_decap_8 FILLER_18_571 ();
 sg13g2_decap_8 FILLER_18_578 ();
 sg13g2_decap_8 FILLER_18_585 ();
 sg13g2_decap_8 FILLER_18_592 ();
 sg13g2_decap_8 FILLER_18_599 ();
 sg13g2_decap_8 FILLER_18_606 ();
 sg13g2_decap_8 FILLER_18_613 ();
 sg13g2_decap_8 FILLER_18_620 ();
 sg13g2_decap_8 FILLER_18_627 ();
 sg13g2_decap_8 FILLER_18_634 ();
 sg13g2_decap_8 FILLER_18_641 ();
 sg13g2_decap_8 FILLER_18_648 ();
 sg13g2_decap_8 FILLER_18_655 ();
 sg13g2_decap_8 FILLER_18_662 ();
 sg13g2_decap_8 FILLER_18_669 ();
 sg13g2_decap_8 FILLER_18_676 ();
 sg13g2_decap_8 FILLER_18_683 ();
 sg13g2_decap_8 FILLER_18_690 ();
 sg13g2_decap_8 FILLER_18_697 ();
 sg13g2_decap_8 FILLER_18_704 ();
 sg13g2_decap_8 FILLER_18_711 ();
 sg13g2_decap_8 FILLER_18_718 ();
 sg13g2_decap_8 FILLER_18_725 ();
 sg13g2_decap_8 FILLER_18_732 ();
 sg13g2_decap_8 FILLER_18_739 ();
 sg13g2_decap_8 FILLER_18_746 ();
 sg13g2_decap_8 FILLER_18_753 ();
 sg13g2_decap_8 FILLER_18_760 ();
 sg13g2_decap_8 FILLER_18_767 ();
 sg13g2_decap_8 FILLER_18_774 ();
 sg13g2_decap_8 FILLER_18_781 ();
 sg13g2_decap_8 FILLER_18_788 ();
 sg13g2_decap_8 FILLER_18_795 ();
 sg13g2_decap_8 FILLER_18_802 ();
 sg13g2_decap_8 FILLER_18_809 ();
 sg13g2_decap_8 FILLER_18_816 ();
 sg13g2_decap_8 FILLER_18_823 ();
 sg13g2_decap_8 FILLER_18_830 ();
 sg13g2_decap_8 FILLER_18_837 ();
 sg13g2_decap_8 FILLER_18_844 ();
 sg13g2_decap_8 FILLER_18_851 ();
 sg13g2_decap_8 FILLER_18_858 ();
 sg13g2_decap_8 FILLER_18_865 ();
 sg13g2_decap_8 FILLER_18_872 ();
 sg13g2_decap_8 FILLER_18_879 ();
 sg13g2_decap_8 FILLER_18_886 ();
 sg13g2_decap_8 FILLER_18_893 ();
 sg13g2_decap_8 FILLER_18_900 ();
 sg13g2_decap_8 FILLER_18_907 ();
 sg13g2_decap_8 FILLER_18_914 ();
 sg13g2_decap_8 FILLER_18_921 ();
 sg13g2_decap_8 FILLER_18_928 ();
 sg13g2_decap_8 FILLER_18_935 ();
 sg13g2_decap_8 FILLER_18_942 ();
 sg13g2_decap_8 FILLER_18_949 ();
 sg13g2_decap_8 FILLER_18_956 ();
 sg13g2_decap_8 FILLER_18_963 ();
 sg13g2_decap_8 FILLER_18_970 ();
 sg13g2_decap_8 FILLER_18_977 ();
 sg13g2_decap_8 FILLER_18_984 ();
 sg13g2_decap_8 FILLER_18_991 ();
 sg13g2_decap_8 FILLER_18_998 ();
 sg13g2_decap_8 FILLER_18_1005 ();
 sg13g2_decap_8 FILLER_18_1012 ();
 sg13g2_decap_8 FILLER_18_1019 ();
 sg13g2_fill_2 FILLER_18_1026 ();
 sg13g2_fill_1 FILLER_18_1028 ();
 sg13g2_decap_8 FILLER_19_4 ();
 sg13g2_decap_8 FILLER_19_11 ();
 sg13g2_decap_8 FILLER_19_18 ();
 sg13g2_decap_8 FILLER_19_25 ();
 sg13g2_decap_8 FILLER_19_32 ();
 sg13g2_decap_8 FILLER_19_39 ();
 sg13g2_decap_8 FILLER_19_46 ();
 sg13g2_decap_8 FILLER_19_53 ();
 sg13g2_decap_8 FILLER_19_60 ();
 sg13g2_decap_8 FILLER_19_67 ();
 sg13g2_decap_8 FILLER_19_74 ();
 sg13g2_decap_8 FILLER_19_81 ();
 sg13g2_decap_8 FILLER_19_88 ();
 sg13g2_decap_8 FILLER_19_95 ();
 sg13g2_decap_8 FILLER_19_102 ();
 sg13g2_decap_8 FILLER_19_109 ();
 sg13g2_decap_8 FILLER_19_116 ();
 sg13g2_decap_8 FILLER_19_123 ();
 sg13g2_decap_8 FILLER_19_130 ();
 sg13g2_decap_8 FILLER_19_137 ();
 sg13g2_decap_8 FILLER_19_144 ();
 sg13g2_fill_2 FILLER_19_151 ();
 sg13g2_fill_1 FILLER_19_153 ();
 sg13g2_fill_2 FILLER_19_181 ();
 sg13g2_decap_8 FILLER_19_192 ();
 sg13g2_decap_8 FILLER_19_199 ();
 sg13g2_decap_8 FILLER_19_206 ();
 sg13g2_decap_8 FILLER_19_213 ();
 sg13g2_decap_8 FILLER_19_220 ();
 sg13g2_decap_8 FILLER_19_227 ();
 sg13g2_decap_8 FILLER_19_234 ();
 sg13g2_decap_8 FILLER_19_241 ();
 sg13g2_decap_8 FILLER_19_248 ();
 sg13g2_decap_8 FILLER_19_255 ();
 sg13g2_decap_8 FILLER_19_262 ();
 sg13g2_decap_8 FILLER_19_269 ();
 sg13g2_decap_8 FILLER_19_276 ();
 sg13g2_fill_1 FILLER_19_283 ();
 sg13g2_decap_8 FILLER_19_290 ();
 sg13g2_decap_8 FILLER_19_297 ();
 sg13g2_decap_8 FILLER_19_304 ();
 sg13g2_decap_8 FILLER_19_311 ();
 sg13g2_decap_8 FILLER_19_318 ();
 sg13g2_decap_8 FILLER_19_325 ();
 sg13g2_decap_8 FILLER_19_332 ();
 sg13g2_decap_8 FILLER_19_339 ();
 sg13g2_decap_8 FILLER_19_346 ();
 sg13g2_decap_8 FILLER_19_353 ();
 sg13g2_decap_8 FILLER_19_360 ();
 sg13g2_decap_8 FILLER_19_367 ();
 sg13g2_decap_8 FILLER_19_374 ();
 sg13g2_decap_4 FILLER_19_381 ();
 sg13g2_decap_8 FILLER_19_412 ();
 sg13g2_decap_8 FILLER_19_419 ();
 sg13g2_decap_8 FILLER_19_426 ();
 sg13g2_decap_8 FILLER_19_433 ();
 sg13g2_decap_8 FILLER_19_440 ();
 sg13g2_decap_8 FILLER_19_447 ();
 sg13g2_decap_8 FILLER_19_454 ();
 sg13g2_decap_8 FILLER_19_461 ();
 sg13g2_decap_8 FILLER_19_468 ();
 sg13g2_decap_8 FILLER_19_475 ();
 sg13g2_decap_8 FILLER_19_482 ();
 sg13g2_decap_8 FILLER_19_489 ();
 sg13g2_decap_8 FILLER_19_496 ();
 sg13g2_decap_8 FILLER_19_503 ();
 sg13g2_decap_8 FILLER_19_510 ();
 sg13g2_decap_8 FILLER_19_517 ();
 sg13g2_decap_8 FILLER_19_524 ();
 sg13g2_decap_8 FILLER_19_531 ();
 sg13g2_decap_8 FILLER_19_538 ();
 sg13g2_decap_8 FILLER_19_545 ();
 sg13g2_decap_8 FILLER_19_552 ();
 sg13g2_decap_8 FILLER_19_559 ();
 sg13g2_decap_8 FILLER_19_566 ();
 sg13g2_decap_8 FILLER_19_573 ();
 sg13g2_decap_8 FILLER_19_580 ();
 sg13g2_decap_8 FILLER_19_587 ();
 sg13g2_decap_8 FILLER_19_594 ();
 sg13g2_decap_8 FILLER_19_601 ();
 sg13g2_decap_8 FILLER_19_608 ();
 sg13g2_decap_8 FILLER_19_615 ();
 sg13g2_decap_8 FILLER_19_622 ();
 sg13g2_decap_8 FILLER_19_629 ();
 sg13g2_decap_8 FILLER_19_636 ();
 sg13g2_decap_8 FILLER_19_643 ();
 sg13g2_decap_8 FILLER_19_650 ();
 sg13g2_decap_8 FILLER_19_657 ();
 sg13g2_decap_8 FILLER_19_664 ();
 sg13g2_decap_8 FILLER_19_671 ();
 sg13g2_decap_8 FILLER_19_678 ();
 sg13g2_decap_8 FILLER_19_685 ();
 sg13g2_decap_8 FILLER_19_692 ();
 sg13g2_decap_8 FILLER_19_699 ();
 sg13g2_decap_8 FILLER_19_706 ();
 sg13g2_decap_8 FILLER_19_713 ();
 sg13g2_decap_8 FILLER_19_720 ();
 sg13g2_decap_8 FILLER_19_727 ();
 sg13g2_decap_8 FILLER_19_734 ();
 sg13g2_decap_8 FILLER_19_741 ();
 sg13g2_decap_8 FILLER_19_748 ();
 sg13g2_decap_8 FILLER_19_755 ();
 sg13g2_decap_8 FILLER_19_762 ();
 sg13g2_decap_8 FILLER_19_769 ();
 sg13g2_decap_8 FILLER_19_776 ();
 sg13g2_decap_8 FILLER_19_783 ();
 sg13g2_decap_8 FILLER_19_790 ();
 sg13g2_decap_8 FILLER_19_797 ();
 sg13g2_decap_8 FILLER_19_804 ();
 sg13g2_decap_8 FILLER_19_811 ();
 sg13g2_decap_8 FILLER_19_818 ();
 sg13g2_decap_8 FILLER_19_825 ();
 sg13g2_decap_8 FILLER_19_832 ();
 sg13g2_decap_8 FILLER_19_839 ();
 sg13g2_decap_8 FILLER_19_846 ();
 sg13g2_decap_8 FILLER_19_853 ();
 sg13g2_decap_8 FILLER_19_860 ();
 sg13g2_decap_8 FILLER_19_867 ();
 sg13g2_decap_8 FILLER_19_874 ();
 sg13g2_decap_8 FILLER_19_881 ();
 sg13g2_decap_8 FILLER_19_888 ();
 sg13g2_decap_8 FILLER_19_895 ();
 sg13g2_decap_8 FILLER_19_902 ();
 sg13g2_decap_8 FILLER_19_909 ();
 sg13g2_decap_8 FILLER_19_916 ();
 sg13g2_decap_8 FILLER_19_923 ();
 sg13g2_decap_8 FILLER_19_930 ();
 sg13g2_decap_8 FILLER_19_937 ();
 sg13g2_decap_8 FILLER_19_944 ();
 sg13g2_decap_8 FILLER_19_951 ();
 sg13g2_decap_8 FILLER_19_958 ();
 sg13g2_decap_8 FILLER_19_965 ();
 sg13g2_decap_8 FILLER_19_972 ();
 sg13g2_decap_8 FILLER_19_979 ();
 sg13g2_decap_8 FILLER_19_986 ();
 sg13g2_decap_8 FILLER_19_993 ();
 sg13g2_decap_8 FILLER_19_1000 ();
 sg13g2_decap_8 FILLER_19_1007 ();
 sg13g2_decap_8 FILLER_19_1014 ();
 sg13g2_decap_8 FILLER_19_1021 ();
 sg13g2_fill_1 FILLER_19_1028 ();
 sg13g2_decap_8 FILLER_20_4 ();
 sg13g2_decap_8 FILLER_20_11 ();
 sg13g2_decap_8 FILLER_20_18 ();
 sg13g2_decap_8 FILLER_20_25 ();
 sg13g2_decap_8 FILLER_20_32 ();
 sg13g2_decap_8 FILLER_20_39 ();
 sg13g2_decap_8 FILLER_20_46 ();
 sg13g2_decap_8 FILLER_20_53 ();
 sg13g2_decap_8 FILLER_20_60 ();
 sg13g2_decap_8 FILLER_20_67 ();
 sg13g2_decap_8 FILLER_20_74 ();
 sg13g2_decap_8 FILLER_20_81 ();
 sg13g2_decap_8 FILLER_20_88 ();
 sg13g2_decap_8 FILLER_20_95 ();
 sg13g2_decap_8 FILLER_20_102 ();
 sg13g2_decap_8 FILLER_20_109 ();
 sg13g2_decap_8 FILLER_20_116 ();
 sg13g2_decap_8 FILLER_20_123 ();
 sg13g2_decap_8 FILLER_20_130 ();
 sg13g2_decap_8 FILLER_20_137 ();
 sg13g2_decap_8 FILLER_20_144 ();
 sg13g2_decap_8 FILLER_20_151 ();
 sg13g2_decap_8 FILLER_20_158 ();
 sg13g2_decap_8 FILLER_20_165 ();
 sg13g2_decap_8 FILLER_20_172 ();
 sg13g2_decap_8 FILLER_20_179 ();
 sg13g2_decap_8 FILLER_20_186 ();
 sg13g2_decap_8 FILLER_20_193 ();
 sg13g2_decap_8 FILLER_20_200 ();
 sg13g2_decap_8 FILLER_20_207 ();
 sg13g2_decap_8 FILLER_20_214 ();
 sg13g2_decap_8 FILLER_20_221 ();
 sg13g2_decap_8 FILLER_20_228 ();
 sg13g2_decap_8 FILLER_20_235 ();
 sg13g2_decap_8 FILLER_20_242 ();
 sg13g2_decap_8 FILLER_20_249 ();
 sg13g2_decap_8 FILLER_20_256 ();
 sg13g2_decap_8 FILLER_20_263 ();
 sg13g2_decap_8 FILLER_20_270 ();
 sg13g2_decap_8 FILLER_20_277 ();
 sg13g2_decap_8 FILLER_20_284 ();
 sg13g2_decap_8 FILLER_20_291 ();
 sg13g2_decap_8 FILLER_20_298 ();
 sg13g2_decap_8 FILLER_20_305 ();
 sg13g2_decap_8 FILLER_20_312 ();
 sg13g2_decap_8 FILLER_20_319 ();
 sg13g2_decap_8 FILLER_20_326 ();
 sg13g2_decap_8 FILLER_20_333 ();
 sg13g2_decap_4 FILLER_20_340 ();
 sg13g2_fill_1 FILLER_20_344 ();
 sg13g2_decap_8 FILLER_20_351 ();
 sg13g2_decap_8 FILLER_20_358 ();
 sg13g2_decap_8 FILLER_20_365 ();
 sg13g2_decap_8 FILLER_20_372 ();
 sg13g2_decap_8 FILLER_20_384 ();
 sg13g2_decap_4 FILLER_20_391 ();
 sg13g2_decap_8 FILLER_20_404 ();
 sg13g2_decap_8 FILLER_20_411 ();
 sg13g2_decap_8 FILLER_20_418 ();
 sg13g2_decap_8 FILLER_20_425 ();
 sg13g2_decap_8 FILLER_20_432 ();
 sg13g2_decap_8 FILLER_20_439 ();
 sg13g2_decap_8 FILLER_20_446 ();
 sg13g2_decap_8 FILLER_20_453 ();
 sg13g2_decap_8 FILLER_20_460 ();
 sg13g2_decap_8 FILLER_20_467 ();
 sg13g2_decap_8 FILLER_20_474 ();
 sg13g2_decap_8 FILLER_20_481 ();
 sg13g2_decap_8 FILLER_20_488 ();
 sg13g2_decap_8 FILLER_20_495 ();
 sg13g2_decap_8 FILLER_20_502 ();
 sg13g2_decap_8 FILLER_20_509 ();
 sg13g2_decap_8 FILLER_20_516 ();
 sg13g2_decap_8 FILLER_20_523 ();
 sg13g2_decap_8 FILLER_20_530 ();
 sg13g2_decap_8 FILLER_20_537 ();
 sg13g2_decap_8 FILLER_20_544 ();
 sg13g2_decap_8 FILLER_20_551 ();
 sg13g2_decap_8 FILLER_20_558 ();
 sg13g2_decap_8 FILLER_20_565 ();
 sg13g2_decap_8 FILLER_20_572 ();
 sg13g2_decap_8 FILLER_20_579 ();
 sg13g2_decap_8 FILLER_20_586 ();
 sg13g2_decap_8 FILLER_20_593 ();
 sg13g2_decap_8 FILLER_20_600 ();
 sg13g2_decap_8 FILLER_20_607 ();
 sg13g2_decap_8 FILLER_20_614 ();
 sg13g2_decap_8 FILLER_20_621 ();
 sg13g2_decap_8 FILLER_20_628 ();
 sg13g2_decap_8 FILLER_20_635 ();
 sg13g2_decap_8 FILLER_20_642 ();
 sg13g2_decap_8 FILLER_20_649 ();
 sg13g2_decap_8 FILLER_20_656 ();
 sg13g2_decap_8 FILLER_20_663 ();
 sg13g2_decap_8 FILLER_20_670 ();
 sg13g2_decap_8 FILLER_20_677 ();
 sg13g2_decap_8 FILLER_20_684 ();
 sg13g2_decap_8 FILLER_20_691 ();
 sg13g2_decap_8 FILLER_20_698 ();
 sg13g2_decap_8 FILLER_20_705 ();
 sg13g2_decap_8 FILLER_20_712 ();
 sg13g2_decap_8 FILLER_20_719 ();
 sg13g2_decap_8 FILLER_20_726 ();
 sg13g2_decap_8 FILLER_20_733 ();
 sg13g2_decap_8 FILLER_20_740 ();
 sg13g2_decap_8 FILLER_20_747 ();
 sg13g2_decap_8 FILLER_20_754 ();
 sg13g2_decap_8 FILLER_20_761 ();
 sg13g2_decap_8 FILLER_20_768 ();
 sg13g2_decap_8 FILLER_20_775 ();
 sg13g2_decap_8 FILLER_20_782 ();
 sg13g2_decap_8 FILLER_20_789 ();
 sg13g2_decap_8 FILLER_20_796 ();
 sg13g2_decap_8 FILLER_20_803 ();
 sg13g2_decap_8 FILLER_20_810 ();
 sg13g2_decap_8 FILLER_20_817 ();
 sg13g2_decap_8 FILLER_20_824 ();
 sg13g2_decap_8 FILLER_20_831 ();
 sg13g2_decap_8 FILLER_20_838 ();
 sg13g2_decap_8 FILLER_20_845 ();
 sg13g2_decap_8 FILLER_20_852 ();
 sg13g2_decap_8 FILLER_20_859 ();
 sg13g2_decap_8 FILLER_20_866 ();
 sg13g2_decap_8 FILLER_20_873 ();
 sg13g2_decap_8 FILLER_20_880 ();
 sg13g2_decap_8 FILLER_20_887 ();
 sg13g2_decap_8 FILLER_20_894 ();
 sg13g2_decap_8 FILLER_20_901 ();
 sg13g2_decap_8 FILLER_20_908 ();
 sg13g2_decap_8 FILLER_20_915 ();
 sg13g2_decap_8 FILLER_20_922 ();
 sg13g2_decap_8 FILLER_20_929 ();
 sg13g2_decap_8 FILLER_20_936 ();
 sg13g2_decap_8 FILLER_20_943 ();
 sg13g2_decap_8 FILLER_20_950 ();
 sg13g2_decap_8 FILLER_20_957 ();
 sg13g2_decap_8 FILLER_20_964 ();
 sg13g2_decap_8 FILLER_20_971 ();
 sg13g2_decap_8 FILLER_20_978 ();
 sg13g2_decap_8 FILLER_20_985 ();
 sg13g2_decap_8 FILLER_20_992 ();
 sg13g2_decap_8 FILLER_20_999 ();
 sg13g2_decap_8 FILLER_20_1006 ();
 sg13g2_decap_8 FILLER_20_1013 ();
 sg13g2_decap_8 FILLER_20_1020 ();
 sg13g2_fill_2 FILLER_20_1027 ();
 sg13g2_decap_8 FILLER_21_4 ();
 sg13g2_decap_8 FILLER_21_11 ();
 sg13g2_decap_8 FILLER_21_18 ();
 sg13g2_decap_8 FILLER_21_25 ();
 sg13g2_decap_8 FILLER_21_32 ();
 sg13g2_decap_8 FILLER_21_39 ();
 sg13g2_decap_8 FILLER_21_46 ();
 sg13g2_decap_8 FILLER_21_53 ();
 sg13g2_decap_8 FILLER_21_60 ();
 sg13g2_decap_8 FILLER_21_67 ();
 sg13g2_decap_8 FILLER_21_74 ();
 sg13g2_decap_8 FILLER_21_81 ();
 sg13g2_decap_8 FILLER_21_88 ();
 sg13g2_decap_8 FILLER_21_95 ();
 sg13g2_decap_8 FILLER_21_102 ();
 sg13g2_decap_8 FILLER_21_109 ();
 sg13g2_decap_8 FILLER_21_116 ();
 sg13g2_decap_8 FILLER_21_123 ();
 sg13g2_decap_8 FILLER_21_130 ();
 sg13g2_decap_8 FILLER_21_137 ();
 sg13g2_decap_8 FILLER_21_144 ();
 sg13g2_decap_8 FILLER_21_151 ();
 sg13g2_decap_8 FILLER_21_162 ();
 sg13g2_decap_8 FILLER_21_169 ();
 sg13g2_decap_8 FILLER_21_176 ();
 sg13g2_decap_8 FILLER_21_183 ();
 sg13g2_decap_8 FILLER_21_190 ();
 sg13g2_decap_8 FILLER_21_197 ();
 sg13g2_decap_8 FILLER_21_204 ();
 sg13g2_decap_8 FILLER_21_211 ();
 sg13g2_decap_4 FILLER_21_218 ();
 sg13g2_fill_1 FILLER_21_222 ();
 sg13g2_decap_8 FILLER_21_228 ();
 sg13g2_decap_8 FILLER_21_235 ();
 sg13g2_decap_8 FILLER_21_242 ();
 sg13g2_decap_8 FILLER_21_249 ();
 sg13g2_decap_8 FILLER_21_256 ();
 sg13g2_decap_8 FILLER_21_263 ();
 sg13g2_decap_8 FILLER_21_270 ();
 sg13g2_decap_8 FILLER_21_277 ();
 sg13g2_decap_8 FILLER_21_284 ();
 sg13g2_decap_8 FILLER_21_291 ();
 sg13g2_decap_8 FILLER_21_298 ();
 sg13g2_decap_8 FILLER_21_305 ();
 sg13g2_decap_8 FILLER_21_312 ();
 sg13g2_fill_1 FILLER_21_319 ();
 sg13g2_decap_8 FILLER_21_353 ();
 sg13g2_decap_8 FILLER_21_360 ();
 sg13g2_decap_8 FILLER_21_367 ();
 sg13g2_decap_8 FILLER_21_374 ();
 sg13g2_decap_8 FILLER_21_381 ();
 sg13g2_decap_8 FILLER_21_388 ();
 sg13g2_decap_8 FILLER_21_395 ();
 sg13g2_decap_8 FILLER_21_402 ();
 sg13g2_decap_8 FILLER_21_409 ();
 sg13g2_decap_8 FILLER_21_416 ();
 sg13g2_decap_8 FILLER_21_423 ();
 sg13g2_decap_8 FILLER_21_430 ();
 sg13g2_decap_8 FILLER_21_437 ();
 sg13g2_decap_8 FILLER_21_444 ();
 sg13g2_decap_8 FILLER_21_451 ();
 sg13g2_decap_8 FILLER_21_458 ();
 sg13g2_decap_8 FILLER_21_465 ();
 sg13g2_decap_8 FILLER_21_472 ();
 sg13g2_decap_8 FILLER_21_479 ();
 sg13g2_decap_8 FILLER_21_486 ();
 sg13g2_decap_8 FILLER_21_493 ();
 sg13g2_decap_8 FILLER_21_500 ();
 sg13g2_decap_8 FILLER_21_507 ();
 sg13g2_decap_8 FILLER_21_514 ();
 sg13g2_decap_8 FILLER_21_521 ();
 sg13g2_decap_8 FILLER_21_528 ();
 sg13g2_decap_8 FILLER_21_535 ();
 sg13g2_decap_8 FILLER_21_542 ();
 sg13g2_decap_8 FILLER_21_549 ();
 sg13g2_decap_8 FILLER_21_556 ();
 sg13g2_decap_8 FILLER_21_563 ();
 sg13g2_decap_8 FILLER_21_570 ();
 sg13g2_decap_8 FILLER_21_577 ();
 sg13g2_decap_8 FILLER_21_584 ();
 sg13g2_decap_8 FILLER_21_591 ();
 sg13g2_decap_8 FILLER_21_598 ();
 sg13g2_decap_8 FILLER_21_605 ();
 sg13g2_decap_8 FILLER_21_612 ();
 sg13g2_decap_8 FILLER_21_619 ();
 sg13g2_decap_8 FILLER_21_626 ();
 sg13g2_decap_8 FILLER_21_633 ();
 sg13g2_decap_8 FILLER_21_640 ();
 sg13g2_decap_8 FILLER_21_647 ();
 sg13g2_decap_8 FILLER_21_654 ();
 sg13g2_decap_8 FILLER_21_661 ();
 sg13g2_decap_8 FILLER_21_668 ();
 sg13g2_decap_8 FILLER_21_675 ();
 sg13g2_decap_8 FILLER_21_682 ();
 sg13g2_decap_8 FILLER_21_689 ();
 sg13g2_decap_8 FILLER_21_696 ();
 sg13g2_decap_8 FILLER_21_703 ();
 sg13g2_decap_8 FILLER_21_710 ();
 sg13g2_decap_8 FILLER_21_717 ();
 sg13g2_decap_8 FILLER_21_724 ();
 sg13g2_decap_8 FILLER_21_731 ();
 sg13g2_decap_8 FILLER_21_738 ();
 sg13g2_decap_8 FILLER_21_745 ();
 sg13g2_decap_8 FILLER_21_752 ();
 sg13g2_decap_8 FILLER_21_759 ();
 sg13g2_decap_8 FILLER_21_766 ();
 sg13g2_decap_8 FILLER_21_773 ();
 sg13g2_decap_8 FILLER_21_780 ();
 sg13g2_decap_8 FILLER_21_787 ();
 sg13g2_decap_8 FILLER_21_794 ();
 sg13g2_decap_8 FILLER_21_801 ();
 sg13g2_decap_8 FILLER_21_808 ();
 sg13g2_decap_8 FILLER_21_815 ();
 sg13g2_decap_8 FILLER_21_822 ();
 sg13g2_decap_8 FILLER_21_829 ();
 sg13g2_decap_8 FILLER_21_836 ();
 sg13g2_decap_8 FILLER_21_843 ();
 sg13g2_decap_8 FILLER_21_850 ();
 sg13g2_decap_8 FILLER_21_857 ();
 sg13g2_decap_8 FILLER_21_864 ();
 sg13g2_decap_8 FILLER_21_871 ();
 sg13g2_decap_8 FILLER_21_878 ();
 sg13g2_decap_8 FILLER_21_885 ();
 sg13g2_decap_8 FILLER_21_892 ();
 sg13g2_decap_8 FILLER_21_899 ();
 sg13g2_decap_8 FILLER_21_906 ();
 sg13g2_decap_8 FILLER_21_913 ();
 sg13g2_decap_8 FILLER_21_920 ();
 sg13g2_decap_8 FILLER_21_927 ();
 sg13g2_decap_8 FILLER_21_934 ();
 sg13g2_decap_8 FILLER_21_941 ();
 sg13g2_decap_8 FILLER_21_948 ();
 sg13g2_decap_8 FILLER_21_955 ();
 sg13g2_decap_8 FILLER_21_962 ();
 sg13g2_decap_8 FILLER_21_969 ();
 sg13g2_decap_8 FILLER_21_976 ();
 sg13g2_decap_8 FILLER_21_983 ();
 sg13g2_decap_8 FILLER_21_990 ();
 sg13g2_decap_8 FILLER_21_997 ();
 sg13g2_decap_8 FILLER_21_1004 ();
 sg13g2_decap_8 FILLER_21_1011 ();
 sg13g2_decap_8 FILLER_21_1018 ();
 sg13g2_decap_4 FILLER_21_1025 ();
 sg13g2_decap_8 FILLER_22_4 ();
 sg13g2_decap_8 FILLER_22_11 ();
 sg13g2_decap_8 FILLER_22_18 ();
 sg13g2_decap_8 FILLER_22_25 ();
 sg13g2_decap_8 FILLER_22_32 ();
 sg13g2_decap_8 FILLER_22_39 ();
 sg13g2_decap_8 FILLER_22_46 ();
 sg13g2_decap_8 FILLER_22_53 ();
 sg13g2_decap_8 FILLER_22_60 ();
 sg13g2_decap_8 FILLER_22_67 ();
 sg13g2_decap_8 FILLER_22_74 ();
 sg13g2_decap_8 FILLER_22_81 ();
 sg13g2_decap_8 FILLER_22_88 ();
 sg13g2_decap_8 FILLER_22_95 ();
 sg13g2_decap_8 FILLER_22_102 ();
 sg13g2_decap_8 FILLER_22_109 ();
 sg13g2_decap_8 FILLER_22_116 ();
 sg13g2_decap_8 FILLER_22_123 ();
 sg13g2_decap_8 FILLER_22_130 ();
 sg13g2_decap_8 FILLER_22_137 ();
 sg13g2_decap_8 FILLER_22_144 ();
 sg13g2_decap_8 FILLER_22_151 ();
 sg13g2_decap_8 FILLER_22_166 ();
 sg13g2_decap_8 FILLER_22_173 ();
 sg13g2_decap_8 FILLER_22_180 ();
 sg13g2_decap_8 FILLER_22_187 ();
 sg13g2_decap_8 FILLER_22_194 ();
 sg13g2_decap_8 FILLER_22_201 ();
 sg13g2_decap_8 FILLER_22_208 ();
 sg13g2_fill_2 FILLER_22_218 ();
 sg13g2_fill_1 FILLER_22_223 ();
 sg13g2_decap_8 FILLER_22_233 ();
 sg13g2_decap_8 FILLER_22_240 ();
 sg13g2_decap_8 FILLER_22_247 ();
 sg13g2_decap_8 FILLER_22_254 ();
 sg13g2_decap_8 FILLER_22_261 ();
 sg13g2_decap_4 FILLER_22_268 ();
 sg13g2_decap_8 FILLER_22_299 ();
 sg13g2_decap_8 FILLER_22_306 ();
 sg13g2_decap_8 FILLER_22_313 ();
 sg13g2_decap_8 FILLER_22_320 ();
 sg13g2_decap_8 FILLER_22_327 ();
 sg13g2_decap_8 FILLER_22_334 ();
 sg13g2_fill_2 FILLER_22_341 ();
 sg13g2_fill_1 FILLER_22_343 ();
 sg13g2_decap_8 FILLER_22_348 ();
 sg13g2_decap_8 FILLER_22_355 ();
 sg13g2_decap_8 FILLER_22_362 ();
 sg13g2_decap_8 FILLER_22_369 ();
 sg13g2_decap_8 FILLER_22_376 ();
 sg13g2_decap_4 FILLER_22_383 ();
 sg13g2_fill_1 FILLER_22_387 ();
 sg13g2_decap_8 FILLER_22_401 ();
 sg13g2_decap_8 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_22_415 ();
 sg13g2_decap_8 FILLER_22_422 ();
 sg13g2_decap_8 FILLER_22_429 ();
 sg13g2_decap_8 FILLER_22_436 ();
 sg13g2_decap_8 FILLER_22_443 ();
 sg13g2_decap_8 FILLER_22_450 ();
 sg13g2_decap_8 FILLER_22_457 ();
 sg13g2_decap_8 FILLER_22_464 ();
 sg13g2_decap_8 FILLER_22_471 ();
 sg13g2_decap_8 FILLER_22_478 ();
 sg13g2_decap_8 FILLER_22_485 ();
 sg13g2_decap_8 FILLER_22_492 ();
 sg13g2_decap_8 FILLER_22_499 ();
 sg13g2_decap_8 FILLER_22_506 ();
 sg13g2_decap_8 FILLER_22_513 ();
 sg13g2_decap_8 FILLER_22_520 ();
 sg13g2_decap_8 FILLER_22_527 ();
 sg13g2_decap_8 FILLER_22_534 ();
 sg13g2_decap_8 FILLER_22_541 ();
 sg13g2_decap_8 FILLER_22_548 ();
 sg13g2_decap_8 FILLER_22_555 ();
 sg13g2_decap_8 FILLER_22_562 ();
 sg13g2_decap_8 FILLER_22_569 ();
 sg13g2_decap_8 FILLER_22_576 ();
 sg13g2_decap_8 FILLER_22_583 ();
 sg13g2_decap_8 FILLER_22_590 ();
 sg13g2_decap_8 FILLER_22_597 ();
 sg13g2_decap_8 FILLER_22_604 ();
 sg13g2_decap_8 FILLER_22_611 ();
 sg13g2_decap_8 FILLER_22_618 ();
 sg13g2_decap_8 FILLER_22_625 ();
 sg13g2_decap_8 FILLER_22_632 ();
 sg13g2_decap_8 FILLER_22_639 ();
 sg13g2_decap_8 FILLER_22_646 ();
 sg13g2_decap_8 FILLER_22_653 ();
 sg13g2_decap_8 FILLER_22_660 ();
 sg13g2_decap_8 FILLER_22_667 ();
 sg13g2_decap_8 FILLER_22_674 ();
 sg13g2_decap_8 FILLER_22_681 ();
 sg13g2_decap_8 FILLER_22_688 ();
 sg13g2_decap_8 FILLER_22_695 ();
 sg13g2_decap_8 FILLER_22_702 ();
 sg13g2_decap_8 FILLER_22_709 ();
 sg13g2_decap_8 FILLER_22_716 ();
 sg13g2_decap_8 FILLER_22_723 ();
 sg13g2_decap_8 FILLER_22_730 ();
 sg13g2_decap_8 FILLER_22_737 ();
 sg13g2_decap_8 FILLER_22_744 ();
 sg13g2_decap_8 FILLER_22_751 ();
 sg13g2_decap_8 FILLER_22_758 ();
 sg13g2_decap_8 FILLER_22_765 ();
 sg13g2_decap_8 FILLER_22_772 ();
 sg13g2_decap_8 FILLER_22_779 ();
 sg13g2_decap_8 FILLER_22_786 ();
 sg13g2_decap_8 FILLER_22_793 ();
 sg13g2_decap_8 FILLER_22_800 ();
 sg13g2_decap_8 FILLER_22_807 ();
 sg13g2_decap_8 FILLER_22_814 ();
 sg13g2_decap_8 FILLER_22_821 ();
 sg13g2_decap_8 FILLER_22_828 ();
 sg13g2_decap_8 FILLER_22_835 ();
 sg13g2_decap_8 FILLER_22_842 ();
 sg13g2_decap_8 FILLER_22_849 ();
 sg13g2_decap_8 FILLER_22_856 ();
 sg13g2_decap_8 FILLER_22_863 ();
 sg13g2_decap_8 FILLER_22_870 ();
 sg13g2_decap_8 FILLER_22_877 ();
 sg13g2_decap_8 FILLER_22_884 ();
 sg13g2_decap_8 FILLER_22_891 ();
 sg13g2_decap_8 FILLER_22_898 ();
 sg13g2_decap_8 FILLER_22_905 ();
 sg13g2_decap_8 FILLER_22_912 ();
 sg13g2_decap_8 FILLER_22_919 ();
 sg13g2_decap_8 FILLER_22_926 ();
 sg13g2_decap_8 FILLER_22_933 ();
 sg13g2_decap_8 FILLER_22_940 ();
 sg13g2_decap_8 FILLER_22_947 ();
 sg13g2_decap_8 FILLER_22_954 ();
 sg13g2_decap_8 FILLER_22_961 ();
 sg13g2_decap_8 FILLER_22_968 ();
 sg13g2_decap_8 FILLER_22_975 ();
 sg13g2_decap_8 FILLER_22_982 ();
 sg13g2_decap_8 FILLER_22_989 ();
 sg13g2_decap_8 FILLER_22_996 ();
 sg13g2_decap_8 FILLER_22_1003 ();
 sg13g2_decap_8 FILLER_22_1010 ();
 sg13g2_decap_8 FILLER_22_1017 ();
 sg13g2_decap_4 FILLER_22_1024 ();
 sg13g2_fill_1 FILLER_22_1028 ();
 sg13g2_decap_8 FILLER_23_4 ();
 sg13g2_decap_8 FILLER_23_11 ();
 sg13g2_decap_8 FILLER_23_18 ();
 sg13g2_decap_8 FILLER_23_25 ();
 sg13g2_decap_8 FILLER_23_32 ();
 sg13g2_decap_8 FILLER_23_39 ();
 sg13g2_decap_8 FILLER_23_46 ();
 sg13g2_decap_8 FILLER_23_53 ();
 sg13g2_decap_8 FILLER_23_60 ();
 sg13g2_decap_8 FILLER_23_67 ();
 sg13g2_decap_8 FILLER_23_74 ();
 sg13g2_decap_8 FILLER_23_81 ();
 sg13g2_decap_8 FILLER_23_88 ();
 sg13g2_decap_8 FILLER_23_95 ();
 sg13g2_decap_8 FILLER_23_102 ();
 sg13g2_decap_8 FILLER_23_109 ();
 sg13g2_decap_8 FILLER_23_116 ();
 sg13g2_decap_8 FILLER_23_123 ();
 sg13g2_decap_8 FILLER_23_130 ();
 sg13g2_decap_8 FILLER_23_137 ();
 sg13g2_decap_8 FILLER_23_144 ();
 sg13g2_decap_8 FILLER_23_151 ();
 sg13g2_decap_8 FILLER_23_158 ();
 sg13g2_decap_8 FILLER_23_165 ();
 sg13g2_fill_2 FILLER_23_172 ();
 sg13g2_fill_1 FILLER_23_174 ();
 sg13g2_decap_8 FILLER_23_183 ();
 sg13g2_decap_8 FILLER_23_190 ();
 sg13g2_decap_8 FILLER_23_197 ();
 sg13g2_decap_8 FILLER_23_204 ();
 sg13g2_decap_8 FILLER_23_211 ();
 sg13g2_decap_4 FILLER_23_218 ();
 sg13g2_fill_2 FILLER_23_222 ();
 sg13g2_decap_8 FILLER_23_230 ();
 sg13g2_decap_8 FILLER_23_237 ();
 sg13g2_decap_8 FILLER_23_244 ();
 sg13g2_decap_8 FILLER_23_251 ();
 sg13g2_decap_8 FILLER_23_258 ();
 sg13g2_decap_8 FILLER_23_271 ();
 sg13g2_decap_8 FILLER_23_281 ();
 sg13g2_fill_1 FILLER_23_288 ();
 sg13g2_decap_8 FILLER_23_298 ();
 sg13g2_decap_8 FILLER_23_305 ();
 sg13g2_decap_8 FILLER_23_312 ();
 sg13g2_decap_8 FILLER_23_319 ();
 sg13g2_decap_8 FILLER_23_326 ();
 sg13g2_decap_8 FILLER_23_333 ();
 sg13g2_decap_8 FILLER_23_340 ();
 sg13g2_decap_8 FILLER_23_347 ();
 sg13g2_decap_8 FILLER_23_354 ();
 sg13g2_decap_8 FILLER_23_361 ();
 sg13g2_decap_8 FILLER_23_368 ();
 sg13g2_decap_8 FILLER_23_375 ();
 sg13g2_decap_8 FILLER_23_382 ();
 sg13g2_decap_8 FILLER_23_389 ();
 sg13g2_decap_8 FILLER_23_396 ();
 sg13g2_decap_8 FILLER_23_403 ();
 sg13g2_decap_8 FILLER_23_410 ();
 sg13g2_decap_8 FILLER_23_417 ();
 sg13g2_decap_8 FILLER_23_424 ();
 sg13g2_decap_8 FILLER_23_431 ();
 sg13g2_decap_8 FILLER_23_438 ();
 sg13g2_decap_8 FILLER_23_445 ();
 sg13g2_decap_8 FILLER_23_452 ();
 sg13g2_decap_8 FILLER_23_459 ();
 sg13g2_decap_8 FILLER_23_466 ();
 sg13g2_decap_8 FILLER_23_473 ();
 sg13g2_decap_8 FILLER_23_480 ();
 sg13g2_decap_8 FILLER_23_487 ();
 sg13g2_decap_8 FILLER_23_494 ();
 sg13g2_decap_8 FILLER_23_501 ();
 sg13g2_decap_8 FILLER_23_508 ();
 sg13g2_decap_8 FILLER_23_515 ();
 sg13g2_decap_8 FILLER_23_522 ();
 sg13g2_decap_8 FILLER_23_529 ();
 sg13g2_decap_8 FILLER_23_536 ();
 sg13g2_decap_8 FILLER_23_543 ();
 sg13g2_decap_8 FILLER_23_550 ();
 sg13g2_decap_8 FILLER_23_557 ();
 sg13g2_decap_8 FILLER_23_564 ();
 sg13g2_decap_8 FILLER_23_571 ();
 sg13g2_decap_8 FILLER_23_578 ();
 sg13g2_decap_8 FILLER_23_585 ();
 sg13g2_decap_8 FILLER_23_592 ();
 sg13g2_decap_8 FILLER_23_599 ();
 sg13g2_decap_8 FILLER_23_606 ();
 sg13g2_decap_8 FILLER_23_613 ();
 sg13g2_decap_8 FILLER_23_620 ();
 sg13g2_decap_8 FILLER_23_627 ();
 sg13g2_decap_8 FILLER_23_634 ();
 sg13g2_decap_8 FILLER_23_641 ();
 sg13g2_decap_8 FILLER_23_648 ();
 sg13g2_decap_8 FILLER_23_655 ();
 sg13g2_decap_8 FILLER_23_662 ();
 sg13g2_decap_8 FILLER_23_669 ();
 sg13g2_decap_8 FILLER_23_676 ();
 sg13g2_decap_8 FILLER_23_683 ();
 sg13g2_decap_8 FILLER_23_690 ();
 sg13g2_decap_8 FILLER_23_697 ();
 sg13g2_decap_8 FILLER_23_704 ();
 sg13g2_decap_8 FILLER_23_711 ();
 sg13g2_decap_8 FILLER_23_718 ();
 sg13g2_decap_8 FILLER_23_725 ();
 sg13g2_decap_8 FILLER_23_732 ();
 sg13g2_decap_8 FILLER_23_739 ();
 sg13g2_decap_8 FILLER_23_746 ();
 sg13g2_decap_8 FILLER_23_753 ();
 sg13g2_decap_8 FILLER_23_760 ();
 sg13g2_decap_8 FILLER_23_767 ();
 sg13g2_decap_8 FILLER_23_774 ();
 sg13g2_decap_8 FILLER_23_781 ();
 sg13g2_decap_8 FILLER_23_788 ();
 sg13g2_decap_8 FILLER_23_795 ();
 sg13g2_decap_8 FILLER_23_802 ();
 sg13g2_decap_8 FILLER_23_809 ();
 sg13g2_decap_8 FILLER_23_816 ();
 sg13g2_decap_8 FILLER_23_823 ();
 sg13g2_decap_8 FILLER_23_830 ();
 sg13g2_decap_8 FILLER_23_837 ();
 sg13g2_decap_8 FILLER_23_844 ();
 sg13g2_decap_8 FILLER_23_851 ();
 sg13g2_decap_8 FILLER_23_858 ();
 sg13g2_decap_8 FILLER_23_865 ();
 sg13g2_decap_8 FILLER_23_872 ();
 sg13g2_decap_8 FILLER_23_879 ();
 sg13g2_decap_8 FILLER_23_886 ();
 sg13g2_decap_8 FILLER_23_893 ();
 sg13g2_decap_8 FILLER_23_900 ();
 sg13g2_decap_8 FILLER_23_907 ();
 sg13g2_decap_8 FILLER_23_914 ();
 sg13g2_decap_8 FILLER_23_921 ();
 sg13g2_decap_8 FILLER_23_928 ();
 sg13g2_decap_8 FILLER_23_935 ();
 sg13g2_decap_8 FILLER_23_942 ();
 sg13g2_decap_8 FILLER_23_949 ();
 sg13g2_decap_8 FILLER_23_956 ();
 sg13g2_decap_8 FILLER_23_963 ();
 sg13g2_decap_8 FILLER_23_970 ();
 sg13g2_decap_8 FILLER_23_977 ();
 sg13g2_decap_8 FILLER_23_984 ();
 sg13g2_decap_8 FILLER_23_991 ();
 sg13g2_decap_8 FILLER_23_998 ();
 sg13g2_decap_8 FILLER_23_1005 ();
 sg13g2_decap_8 FILLER_23_1012 ();
 sg13g2_decap_8 FILLER_23_1019 ();
 sg13g2_fill_2 FILLER_23_1026 ();
 sg13g2_fill_1 FILLER_23_1028 ();
 sg13g2_decap_8 FILLER_24_4 ();
 sg13g2_decap_8 FILLER_24_11 ();
 sg13g2_decap_8 FILLER_24_18 ();
 sg13g2_decap_8 FILLER_24_25 ();
 sg13g2_decap_8 FILLER_24_32 ();
 sg13g2_decap_8 FILLER_24_39 ();
 sg13g2_decap_8 FILLER_24_46 ();
 sg13g2_decap_8 FILLER_24_53 ();
 sg13g2_decap_8 FILLER_24_60 ();
 sg13g2_decap_8 FILLER_24_67 ();
 sg13g2_decap_8 FILLER_24_74 ();
 sg13g2_decap_8 FILLER_24_81 ();
 sg13g2_decap_8 FILLER_24_88 ();
 sg13g2_decap_8 FILLER_24_95 ();
 sg13g2_decap_8 FILLER_24_102 ();
 sg13g2_decap_8 FILLER_24_109 ();
 sg13g2_decap_8 FILLER_24_116 ();
 sg13g2_decap_8 FILLER_24_123 ();
 sg13g2_decap_8 FILLER_24_130 ();
 sg13g2_decap_8 FILLER_24_137 ();
 sg13g2_decap_8 FILLER_24_144 ();
 sg13g2_decap_8 FILLER_24_151 ();
 sg13g2_decap_8 FILLER_24_158 ();
 sg13g2_decap_8 FILLER_24_165 ();
 sg13g2_decap_8 FILLER_24_172 ();
 sg13g2_decap_8 FILLER_24_179 ();
 sg13g2_fill_2 FILLER_24_186 ();
 sg13g2_fill_1 FILLER_24_188 ();
 sg13g2_decap_8 FILLER_24_201 ();
 sg13g2_decap_8 FILLER_24_208 ();
 sg13g2_decap_8 FILLER_24_215 ();
 sg13g2_decap_8 FILLER_24_222 ();
 sg13g2_decap_8 FILLER_24_229 ();
 sg13g2_decap_8 FILLER_24_236 ();
 sg13g2_decap_8 FILLER_24_243 ();
 sg13g2_decap_8 FILLER_24_250 ();
 sg13g2_decap_8 FILLER_24_257 ();
 sg13g2_decap_8 FILLER_24_264 ();
 sg13g2_decap_8 FILLER_24_271 ();
 sg13g2_decap_8 FILLER_24_278 ();
 sg13g2_decap_8 FILLER_24_285 ();
 sg13g2_decap_8 FILLER_24_292 ();
 sg13g2_decap_8 FILLER_24_299 ();
 sg13g2_decap_8 FILLER_24_306 ();
 sg13g2_decap_8 FILLER_24_313 ();
 sg13g2_decap_8 FILLER_24_320 ();
 sg13g2_decap_8 FILLER_24_327 ();
 sg13g2_decap_4 FILLER_24_334 ();
 sg13g2_decap_8 FILLER_24_351 ();
 sg13g2_decap_8 FILLER_24_358 ();
 sg13g2_decap_8 FILLER_24_365 ();
 sg13g2_decap_4 FILLER_24_372 ();
 sg13g2_decap_8 FILLER_24_386 ();
 sg13g2_decap_4 FILLER_24_393 ();
 sg13g2_decap_8 FILLER_24_424 ();
 sg13g2_decap_8 FILLER_24_431 ();
 sg13g2_decap_8 FILLER_24_438 ();
 sg13g2_decap_8 FILLER_24_445 ();
 sg13g2_decap_8 FILLER_24_452 ();
 sg13g2_decap_8 FILLER_24_459 ();
 sg13g2_decap_8 FILLER_24_466 ();
 sg13g2_decap_8 FILLER_24_473 ();
 sg13g2_decap_8 FILLER_24_480 ();
 sg13g2_decap_8 FILLER_24_487 ();
 sg13g2_decap_8 FILLER_24_494 ();
 sg13g2_decap_8 FILLER_24_501 ();
 sg13g2_decap_8 FILLER_24_508 ();
 sg13g2_decap_8 FILLER_24_515 ();
 sg13g2_decap_8 FILLER_24_522 ();
 sg13g2_decap_8 FILLER_24_529 ();
 sg13g2_decap_8 FILLER_24_536 ();
 sg13g2_decap_8 FILLER_24_543 ();
 sg13g2_decap_8 FILLER_24_550 ();
 sg13g2_decap_8 FILLER_24_557 ();
 sg13g2_decap_8 FILLER_24_564 ();
 sg13g2_decap_8 FILLER_24_571 ();
 sg13g2_decap_8 FILLER_24_578 ();
 sg13g2_decap_8 FILLER_24_585 ();
 sg13g2_decap_8 FILLER_24_592 ();
 sg13g2_decap_8 FILLER_24_599 ();
 sg13g2_decap_8 FILLER_24_606 ();
 sg13g2_decap_8 FILLER_24_613 ();
 sg13g2_decap_8 FILLER_24_620 ();
 sg13g2_decap_8 FILLER_24_627 ();
 sg13g2_decap_8 FILLER_24_634 ();
 sg13g2_decap_8 FILLER_24_641 ();
 sg13g2_decap_8 FILLER_24_648 ();
 sg13g2_decap_8 FILLER_24_655 ();
 sg13g2_decap_8 FILLER_24_662 ();
 sg13g2_decap_8 FILLER_24_669 ();
 sg13g2_decap_8 FILLER_24_676 ();
 sg13g2_decap_8 FILLER_24_683 ();
 sg13g2_decap_8 FILLER_24_690 ();
 sg13g2_decap_8 FILLER_24_697 ();
 sg13g2_decap_8 FILLER_24_704 ();
 sg13g2_decap_8 FILLER_24_711 ();
 sg13g2_decap_8 FILLER_24_718 ();
 sg13g2_decap_8 FILLER_24_725 ();
 sg13g2_decap_8 FILLER_24_732 ();
 sg13g2_decap_8 FILLER_24_739 ();
 sg13g2_decap_8 FILLER_24_746 ();
 sg13g2_decap_8 FILLER_24_753 ();
 sg13g2_decap_8 FILLER_24_760 ();
 sg13g2_decap_8 FILLER_24_767 ();
 sg13g2_decap_8 FILLER_24_774 ();
 sg13g2_decap_8 FILLER_24_781 ();
 sg13g2_decap_8 FILLER_24_788 ();
 sg13g2_decap_8 FILLER_24_795 ();
 sg13g2_decap_8 FILLER_24_802 ();
 sg13g2_decap_8 FILLER_24_809 ();
 sg13g2_decap_8 FILLER_24_816 ();
 sg13g2_decap_8 FILLER_24_823 ();
 sg13g2_decap_8 FILLER_24_830 ();
 sg13g2_decap_8 FILLER_24_837 ();
 sg13g2_decap_8 FILLER_24_844 ();
 sg13g2_decap_8 FILLER_24_851 ();
 sg13g2_decap_8 FILLER_24_858 ();
 sg13g2_decap_8 FILLER_24_865 ();
 sg13g2_decap_8 FILLER_24_872 ();
 sg13g2_decap_8 FILLER_24_879 ();
 sg13g2_decap_8 FILLER_24_886 ();
 sg13g2_decap_8 FILLER_24_893 ();
 sg13g2_decap_8 FILLER_24_900 ();
 sg13g2_decap_8 FILLER_24_907 ();
 sg13g2_decap_8 FILLER_24_914 ();
 sg13g2_decap_8 FILLER_24_921 ();
 sg13g2_decap_8 FILLER_24_928 ();
 sg13g2_decap_8 FILLER_24_935 ();
 sg13g2_decap_8 FILLER_24_942 ();
 sg13g2_decap_8 FILLER_24_949 ();
 sg13g2_decap_8 FILLER_24_956 ();
 sg13g2_decap_8 FILLER_24_963 ();
 sg13g2_decap_8 FILLER_24_970 ();
 sg13g2_decap_8 FILLER_24_977 ();
 sg13g2_decap_8 FILLER_24_984 ();
 sg13g2_decap_8 FILLER_24_991 ();
 sg13g2_decap_8 FILLER_24_998 ();
 sg13g2_decap_8 FILLER_24_1005 ();
 sg13g2_decap_8 FILLER_24_1012 ();
 sg13g2_decap_8 FILLER_24_1019 ();
 sg13g2_fill_2 FILLER_24_1026 ();
 sg13g2_fill_1 FILLER_24_1028 ();
 sg13g2_decap_8 FILLER_25_4 ();
 sg13g2_decap_8 FILLER_25_11 ();
 sg13g2_decap_8 FILLER_25_18 ();
 sg13g2_decap_8 FILLER_25_25 ();
 sg13g2_decap_8 FILLER_25_32 ();
 sg13g2_decap_8 FILLER_25_39 ();
 sg13g2_decap_8 FILLER_25_46 ();
 sg13g2_decap_8 FILLER_25_53 ();
 sg13g2_decap_8 FILLER_25_60 ();
 sg13g2_decap_8 FILLER_25_67 ();
 sg13g2_decap_8 FILLER_25_74 ();
 sg13g2_decap_8 FILLER_25_81 ();
 sg13g2_decap_8 FILLER_25_88 ();
 sg13g2_decap_8 FILLER_25_95 ();
 sg13g2_decap_8 FILLER_25_102 ();
 sg13g2_decap_8 FILLER_25_109 ();
 sg13g2_decap_8 FILLER_25_116 ();
 sg13g2_decap_8 FILLER_25_123 ();
 sg13g2_decap_8 FILLER_25_130 ();
 sg13g2_decap_8 FILLER_25_137 ();
 sg13g2_decap_8 FILLER_25_144 ();
 sg13g2_fill_2 FILLER_25_151 ();
 sg13g2_decap_8 FILLER_25_161 ();
 sg13g2_decap_8 FILLER_25_168 ();
 sg13g2_decap_8 FILLER_25_175 ();
 sg13g2_decap_8 FILLER_25_182 ();
 sg13g2_decap_8 FILLER_25_189 ();
 sg13g2_decap_8 FILLER_25_196 ();
 sg13g2_decap_8 FILLER_25_203 ();
 sg13g2_fill_2 FILLER_25_210 ();
 sg13g2_fill_1 FILLER_25_212 ();
 sg13g2_fill_2 FILLER_25_218 ();
 sg13g2_decap_4 FILLER_25_225 ();
 sg13g2_fill_2 FILLER_25_229 ();
 sg13g2_decap_8 FILLER_25_248 ();
 sg13g2_decap_8 FILLER_25_255 ();
 sg13g2_decap_8 FILLER_25_262 ();
 sg13g2_decap_8 FILLER_25_269 ();
 sg13g2_decap_8 FILLER_25_276 ();
 sg13g2_decap_8 FILLER_25_283 ();
 sg13g2_decap_8 FILLER_25_290 ();
 sg13g2_decap_8 FILLER_25_297 ();
 sg13g2_decap_8 FILLER_25_304 ();
 sg13g2_decap_8 FILLER_25_311 ();
 sg13g2_decap_8 FILLER_25_318 ();
 sg13g2_decap_8 FILLER_25_325 ();
 sg13g2_decap_8 FILLER_25_332 ();
 sg13g2_decap_8 FILLER_25_339 ();
 sg13g2_decap_8 FILLER_25_346 ();
 sg13g2_fill_2 FILLER_25_353 ();
 sg13g2_fill_1 FILLER_25_355 ();
 sg13g2_decap_8 FILLER_25_360 ();
 sg13g2_decap_8 FILLER_25_367 ();
 sg13g2_decap_8 FILLER_25_374 ();
 sg13g2_decap_8 FILLER_25_381 ();
 sg13g2_decap_8 FILLER_25_388 ();
 sg13g2_decap_8 FILLER_25_395 ();
 sg13g2_decap_8 FILLER_25_411 ();
 sg13g2_decap_8 FILLER_25_418 ();
 sg13g2_decap_8 FILLER_25_425 ();
 sg13g2_decap_8 FILLER_25_432 ();
 sg13g2_decap_8 FILLER_25_439 ();
 sg13g2_decap_8 FILLER_25_446 ();
 sg13g2_decap_8 FILLER_25_453 ();
 sg13g2_decap_8 FILLER_25_460 ();
 sg13g2_decap_8 FILLER_25_467 ();
 sg13g2_decap_8 FILLER_25_474 ();
 sg13g2_decap_8 FILLER_25_481 ();
 sg13g2_decap_8 FILLER_25_488 ();
 sg13g2_decap_8 FILLER_25_495 ();
 sg13g2_decap_8 FILLER_25_502 ();
 sg13g2_decap_8 FILLER_25_509 ();
 sg13g2_decap_8 FILLER_25_516 ();
 sg13g2_decap_8 FILLER_25_523 ();
 sg13g2_decap_8 FILLER_25_530 ();
 sg13g2_decap_8 FILLER_25_537 ();
 sg13g2_decap_8 FILLER_25_544 ();
 sg13g2_decap_8 FILLER_25_551 ();
 sg13g2_decap_8 FILLER_25_558 ();
 sg13g2_decap_8 FILLER_25_565 ();
 sg13g2_decap_8 FILLER_25_572 ();
 sg13g2_decap_8 FILLER_25_579 ();
 sg13g2_decap_8 FILLER_25_586 ();
 sg13g2_decap_8 FILLER_25_593 ();
 sg13g2_decap_8 FILLER_25_600 ();
 sg13g2_decap_8 FILLER_25_607 ();
 sg13g2_decap_8 FILLER_25_614 ();
 sg13g2_decap_8 FILLER_25_621 ();
 sg13g2_decap_8 FILLER_25_628 ();
 sg13g2_decap_8 FILLER_25_635 ();
 sg13g2_decap_8 FILLER_25_642 ();
 sg13g2_decap_8 FILLER_25_649 ();
 sg13g2_decap_8 FILLER_25_656 ();
 sg13g2_decap_8 FILLER_25_663 ();
 sg13g2_decap_8 FILLER_25_670 ();
 sg13g2_decap_8 FILLER_25_677 ();
 sg13g2_decap_8 FILLER_25_684 ();
 sg13g2_decap_8 FILLER_25_691 ();
 sg13g2_decap_8 FILLER_25_698 ();
 sg13g2_decap_8 FILLER_25_705 ();
 sg13g2_decap_8 FILLER_25_712 ();
 sg13g2_decap_8 FILLER_25_719 ();
 sg13g2_decap_8 FILLER_25_726 ();
 sg13g2_decap_8 FILLER_25_733 ();
 sg13g2_decap_8 FILLER_25_740 ();
 sg13g2_decap_8 FILLER_25_747 ();
 sg13g2_decap_8 FILLER_25_754 ();
 sg13g2_decap_8 FILLER_25_761 ();
 sg13g2_decap_8 FILLER_25_768 ();
 sg13g2_decap_8 FILLER_25_775 ();
 sg13g2_decap_8 FILLER_25_782 ();
 sg13g2_decap_8 FILLER_25_789 ();
 sg13g2_decap_8 FILLER_25_796 ();
 sg13g2_decap_8 FILLER_25_803 ();
 sg13g2_decap_8 FILLER_25_810 ();
 sg13g2_decap_8 FILLER_25_817 ();
 sg13g2_decap_8 FILLER_25_824 ();
 sg13g2_decap_8 FILLER_25_831 ();
 sg13g2_decap_8 FILLER_25_838 ();
 sg13g2_decap_8 FILLER_25_845 ();
 sg13g2_decap_8 FILLER_25_852 ();
 sg13g2_decap_8 FILLER_25_859 ();
 sg13g2_decap_8 FILLER_25_866 ();
 sg13g2_decap_8 FILLER_25_873 ();
 sg13g2_decap_8 FILLER_25_880 ();
 sg13g2_decap_8 FILLER_25_887 ();
 sg13g2_decap_8 FILLER_25_894 ();
 sg13g2_decap_8 FILLER_25_901 ();
 sg13g2_decap_8 FILLER_25_908 ();
 sg13g2_decap_8 FILLER_25_915 ();
 sg13g2_decap_8 FILLER_25_922 ();
 sg13g2_decap_8 FILLER_25_929 ();
 sg13g2_decap_8 FILLER_25_936 ();
 sg13g2_decap_8 FILLER_25_943 ();
 sg13g2_decap_8 FILLER_25_950 ();
 sg13g2_decap_8 FILLER_25_957 ();
 sg13g2_decap_8 FILLER_25_964 ();
 sg13g2_decap_8 FILLER_25_971 ();
 sg13g2_decap_8 FILLER_25_978 ();
 sg13g2_decap_8 FILLER_25_985 ();
 sg13g2_decap_8 FILLER_25_992 ();
 sg13g2_decap_8 FILLER_25_999 ();
 sg13g2_decap_8 FILLER_25_1006 ();
 sg13g2_decap_8 FILLER_25_1013 ();
 sg13g2_decap_8 FILLER_25_1020 ();
 sg13g2_fill_2 FILLER_25_1027 ();
 sg13g2_decap_8 FILLER_26_4 ();
 sg13g2_decap_8 FILLER_26_11 ();
 sg13g2_decap_8 FILLER_26_18 ();
 sg13g2_decap_8 FILLER_26_25 ();
 sg13g2_decap_8 FILLER_26_32 ();
 sg13g2_decap_8 FILLER_26_39 ();
 sg13g2_decap_8 FILLER_26_46 ();
 sg13g2_decap_8 FILLER_26_53 ();
 sg13g2_decap_8 FILLER_26_60 ();
 sg13g2_decap_8 FILLER_26_67 ();
 sg13g2_decap_8 FILLER_26_74 ();
 sg13g2_decap_8 FILLER_26_81 ();
 sg13g2_decap_8 FILLER_26_88 ();
 sg13g2_decap_8 FILLER_26_95 ();
 sg13g2_decap_8 FILLER_26_102 ();
 sg13g2_decap_8 FILLER_26_109 ();
 sg13g2_decap_8 FILLER_26_116 ();
 sg13g2_decap_8 FILLER_26_123 ();
 sg13g2_decap_8 FILLER_26_130 ();
 sg13g2_decap_8 FILLER_26_137 ();
 sg13g2_decap_8 FILLER_26_144 ();
 sg13g2_decap_8 FILLER_26_151 ();
 sg13g2_decap_8 FILLER_26_158 ();
 sg13g2_decap_8 FILLER_26_165 ();
 sg13g2_decap_8 FILLER_26_172 ();
 sg13g2_decap_8 FILLER_26_179 ();
 sg13g2_decap_8 FILLER_26_186 ();
 sg13g2_decap_8 FILLER_26_200 ();
 sg13g2_decap_8 FILLER_26_207 ();
 sg13g2_decap_8 FILLER_26_214 ();
 sg13g2_decap_8 FILLER_26_221 ();
 sg13g2_fill_1 FILLER_26_228 ();
 sg13g2_decap_8 FILLER_26_239 ();
 sg13g2_decap_8 FILLER_26_246 ();
 sg13g2_decap_8 FILLER_26_253 ();
 sg13g2_decap_8 FILLER_26_260 ();
 sg13g2_decap_8 FILLER_26_267 ();
 sg13g2_decap_8 FILLER_26_274 ();
 sg13g2_decap_8 FILLER_26_281 ();
 sg13g2_decap_8 FILLER_26_288 ();
 sg13g2_fill_2 FILLER_26_295 ();
 sg13g2_decap_4 FILLER_26_304 ();
 sg13g2_fill_1 FILLER_26_308 ();
 sg13g2_decap_8 FILLER_26_322 ();
 sg13g2_decap_8 FILLER_26_329 ();
 sg13g2_decap_8 FILLER_26_336 ();
 sg13g2_decap_8 FILLER_26_343 ();
 sg13g2_decap_8 FILLER_26_350 ();
 sg13g2_decap_8 FILLER_26_357 ();
 sg13g2_decap_8 FILLER_26_364 ();
 sg13g2_decap_8 FILLER_26_371 ();
 sg13g2_decap_8 FILLER_26_378 ();
 sg13g2_decap_8 FILLER_26_385 ();
 sg13g2_decap_8 FILLER_26_392 ();
 sg13g2_decap_8 FILLER_26_399 ();
 sg13g2_decap_8 FILLER_26_406 ();
 sg13g2_decap_8 FILLER_26_413 ();
 sg13g2_decap_8 FILLER_26_420 ();
 sg13g2_decap_8 FILLER_26_427 ();
 sg13g2_decap_8 FILLER_26_434 ();
 sg13g2_decap_8 FILLER_26_441 ();
 sg13g2_decap_8 FILLER_26_448 ();
 sg13g2_decap_8 FILLER_26_455 ();
 sg13g2_decap_8 FILLER_26_462 ();
 sg13g2_decap_8 FILLER_26_469 ();
 sg13g2_decap_8 FILLER_26_476 ();
 sg13g2_decap_8 FILLER_26_483 ();
 sg13g2_decap_8 FILLER_26_490 ();
 sg13g2_decap_8 FILLER_26_497 ();
 sg13g2_decap_8 FILLER_26_504 ();
 sg13g2_decap_8 FILLER_26_511 ();
 sg13g2_decap_8 FILLER_26_518 ();
 sg13g2_decap_8 FILLER_26_525 ();
 sg13g2_decap_8 FILLER_26_532 ();
 sg13g2_decap_8 FILLER_26_539 ();
 sg13g2_decap_8 FILLER_26_546 ();
 sg13g2_decap_8 FILLER_26_553 ();
 sg13g2_decap_8 FILLER_26_560 ();
 sg13g2_decap_8 FILLER_26_567 ();
 sg13g2_decap_8 FILLER_26_574 ();
 sg13g2_decap_8 FILLER_26_581 ();
 sg13g2_decap_8 FILLER_26_588 ();
 sg13g2_decap_8 FILLER_26_595 ();
 sg13g2_decap_8 FILLER_26_602 ();
 sg13g2_decap_8 FILLER_26_609 ();
 sg13g2_decap_8 FILLER_26_616 ();
 sg13g2_decap_8 FILLER_26_623 ();
 sg13g2_decap_8 FILLER_26_630 ();
 sg13g2_decap_8 FILLER_26_637 ();
 sg13g2_decap_8 FILLER_26_644 ();
 sg13g2_decap_8 FILLER_26_651 ();
 sg13g2_decap_8 FILLER_26_658 ();
 sg13g2_decap_8 FILLER_26_665 ();
 sg13g2_decap_8 FILLER_26_672 ();
 sg13g2_decap_8 FILLER_26_679 ();
 sg13g2_decap_8 FILLER_26_686 ();
 sg13g2_decap_8 FILLER_26_693 ();
 sg13g2_decap_8 FILLER_26_700 ();
 sg13g2_decap_8 FILLER_26_707 ();
 sg13g2_decap_8 FILLER_26_714 ();
 sg13g2_decap_8 FILLER_26_721 ();
 sg13g2_decap_8 FILLER_26_728 ();
 sg13g2_decap_8 FILLER_26_735 ();
 sg13g2_decap_8 FILLER_26_742 ();
 sg13g2_decap_8 FILLER_26_749 ();
 sg13g2_decap_8 FILLER_26_756 ();
 sg13g2_decap_8 FILLER_26_763 ();
 sg13g2_decap_8 FILLER_26_770 ();
 sg13g2_decap_8 FILLER_26_777 ();
 sg13g2_decap_8 FILLER_26_784 ();
 sg13g2_decap_8 FILLER_26_791 ();
 sg13g2_decap_8 FILLER_26_798 ();
 sg13g2_decap_8 FILLER_26_805 ();
 sg13g2_decap_8 FILLER_26_812 ();
 sg13g2_decap_8 FILLER_26_819 ();
 sg13g2_decap_8 FILLER_26_826 ();
 sg13g2_decap_8 FILLER_26_833 ();
 sg13g2_decap_8 FILLER_26_840 ();
 sg13g2_decap_8 FILLER_26_847 ();
 sg13g2_decap_8 FILLER_26_854 ();
 sg13g2_decap_8 FILLER_26_861 ();
 sg13g2_decap_8 FILLER_26_868 ();
 sg13g2_decap_8 FILLER_26_875 ();
 sg13g2_decap_8 FILLER_26_882 ();
 sg13g2_decap_8 FILLER_26_889 ();
 sg13g2_decap_8 FILLER_26_896 ();
 sg13g2_decap_8 FILLER_26_903 ();
 sg13g2_decap_8 FILLER_26_910 ();
 sg13g2_decap_8 FILLER_26_917 ();
 sg13g2_decap_8 FILLER_26_924 ();
 sg13g2_decap_8 FILLER_26_931 ();
 sg13g2_decap_8 FILLER_26_938 ();
 sg13g2_decap_8 FILLER_26_945 ();
 sg13g2_decap_8 FILLER_26_952 ();
 sg13g2_decap_8 FILLER_26_959 ();
 sg13g2_decap_8 FILLER_26_966 ();
 sg13g2_decap_8 FILLER_26_973 ();
 sg13g2_decap_8 FILLER_26_980 ();
 sg13g2_decap_8 FILLER_26_987 ();
 sg13g2_decap_8 FILLER_26_994 ();
 sg13g2_decap_8 FILLER_26_1001 ();
 sg13g2_decap_8 FILLER_26_1008 ();
 sg13g2_decap_8 FILLER_26_1015 ();
 sg13g2_decap_8 FILLER_26_1022 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_decap_8 FILLER_27_112 ();
 sg13g2_decap_8 FILLER_27_119 ();
 sg13g2_decap_8 FILLER_27_126 ();
 sg13g2_decap_8 FILLER_27_133 ();
 sg13g2_decap_8 FILLER_27_140 ();
 sg13g2_decap_8 FILLER_27_147 ();
 sg13g2_decap_8 FILLER_27_154 ();
 sg13g2_decap_8 FILLER_27_161 ();
 sg13g2_decap_8 FILLER_27_168 ();
 sg13g2_decap_8 FILLER_27_175 ();
 sg13g2_decap_8 FILLER_27_182 ();
 sg13g2_decap_8 FILLER_27_189 ();
 sg13g2_decap_8 FILLER_27_196 ();
 sg13g2_decap_8 FILLER_27_203 ();
 sg13g2_decap_8 FILLER_27_210 ();
 sg13g2_decap_8 FILLER_27_217 ();
 sg13g2_decap_8 FILLER_27_224 ();
 sg13g2_decap_8 FILLER_27_231 ();
 sg13g2_decap_8 FILLER_27_238 ();
 sg13g2_decap_8 FILLER_27_245 ();
 sg13g2_decap_8 FILLER_27_252 ();
 sg13g2_decap_8 FILLER_27_259 ();
 sg13g2_decap_8 FILLER_27_266 ();
 sg13g2_decap_8 FILLER_27_273 ();
 sg13g2_decap_8 FILLER_27_280 ();
 sg13g2_fill_1 FILLER_27_287 ();
 sg13g2_decap_8 FILLER_27_301 ();
 sg13g2_decap_8 FILLER_27_308 ();
 sg13g2_decap_8 FILLER_27_315 ();
 sg13g2_decap_8 FILLER_27_322 ();
 sg13g2_decap_8 FILLER_27_329 ();
 sg13g2_decap_8 FILLER_27_336 ();
 sg13g2_decap_8 FILLER_27_343 ();
 sg13g2_decap_8 FILLER_27_350 ();
 sg13g2_decap_8 FILLER_27_357 ();
 sg13g2_decap_8 FILLER_27_364 ();
 sg13g2_decap_8 FILLER_27_371 ();
 sg13g2_decap_8 FILLER_27_378 ();
 sg13g2_decap_8 FILLER_27_385 ();
 sg13g2_decap_8 FILLER_27_392 ();
 sg13g2_decap_8 FILLER_27_399 ();
 sg13g2_decap_8 FILLER_27_406 ();
 sg13g2_decap_8 FILLER_27_413 ();
 sg13g2_decap_8 FILLER_27_420 ();
 sg13g2_decap_8 FILLER_27_427 ();
 sg13g2_decap_8 FILLER_27_434 ();
 sg13g2_decap_8 FILLER_27_441 ();
 sg13g2_decap_8 FILLER_27_448 ();
 sg13g2_decap_8 FILLER_27_455 ();
 sg13g2_decap_8 FILLER_27_462 ();
 sg13g2_decap_8 FILLER_27_469 ();
 sg13g2_decap_8 FILLER_27_476 ();
 sg13g2_decap_8 FILLER_27_483 ();
 sg13g2_decap_8 FILLER_27_490 ();
 sg13g2_decap_8 FILLER_27_497 ();
 sg13g2_decap_8 FILLER_27_504 ();
 sg13g2_decap_8 FILLER_27_511 ();
 sg13g2_decap_8 FILLER_27_518 ();
 sg13g2_decap_8 FILLER_27_525 ();
 sg13g2_decap_8 FILLER_27_532 ();
 sg13g2_decap_8 FILLER_27_539 ();
 sg13g2_decap_8 FILLER_27_546 ();
 sg13g2_decap_8 FILLER_27_553 ();
 sg13g2_decap_8 FILLER_27_560 ();
 sg13g2_decap_8 FILLER_27_567 ();
 sg13g2_decap_8 FILLER_27_574 ();
 sg13g2_decap_8 FILLER_27_581 ();
 sg13g2_decap_8 FILLER_27_588 ();
 sg13g2_decap_8 FILLER_27_595 ();
 sg13g2_decap_8 FILLER_27_602 ();
 sg13g2_decap_8 FILLER_27_609 ();
 sg13g2_decap_8 FILLER_27_616 ();
 sg13g2_decap_8 FILLER_27_623 ();
 sg13g2_decap_8 FILLER_27_630 ();
 sg13g2_decap_8 FILLER_27_637 ();
 sg13g2_decap_8 FILLER_27_644 ();
 sg13g2_decap_8 FILLER_27_651 ();
 sg13g2_decap_8 FILLER_27_658 ();
 sg13g2_decap_8 FILLER_27_665 ();
 sg13g2_decap_8 FILLER_27_672 ();
 sg13g2_decap_8 FILLER_27_679 ();
 sg13g2_decap_8 FILLER_27_686 ();
 sg13g2_decap_8 FILLER_27_693 ();
 sg13g2_decap_8 FILLER_27_700 ();
 sg13g2_decap_8 FILLER_27_707 ();
 sg13g2_decap_8 FILLER_27_714 ();
 sg13g2_decap_8 FILLER_27_721 ();
 sg13g2_decap_8 FILLER_27_728 ();
 sg13g2_decap_8 FILLER_27_735 ();
 sg13g2_decap_8 FILLER_27_742 ();
 sg13g2_decap_8 FILLER_27_749 ();
 sg13g2_decap_8 FILLER_27_756 ();
 sg13g2_decap_8 FILLER_27_763 ();
 sg13g2_decap_8 FILLER_27_770 ();
 sg13g2_decap_8 FILLER_27_777 ();
 sg13g2_decap_8 FILLER_27_784 ();
 sg13g2_decap_8 FILLER_27_791 ();
 sg13g2_decap_8 FILLER_27_798 ();
 sg13g2_decap_8 FILLER_27_805 ();
 sg13g2_decap_8 FILLER_27_812 ();
 sg13g2_decap_8 FILLER_27_819 ();
 sg13g2_decap_8 FILLER_27_826 ();
 sg13g2_decap_8 FILLER_27_833 ();
 sg13g2_decap_8 FILLER_27_840 ();
 sg13g2_decap_8 FILLER_27_847 ();
 sg13g2_decap_8 FILLER_27_854 ();
 sg13g2_decap_8 FILLER_27_861 ();
 sg13g2_decap_8 FILLER_27_868 ();
 sg13g2_decap_8 FILLER_27_875 ();
 sg13g2_decap_8 FILLER_27_882 ();
 sg13g2_decap_8 FILLER_27_889 ();
 sg13g2_decap_8 FILLER_27_896 ();
 sg13g2_decap_8 FILLER_27_903 ();
 sg13g2_decap_8 FILLER_27_910 ();
 sg13g2_decap_8 FILLER_27_917 ();
 sg13g2_decap_8 FILLER_27_924 ();
 sg13g2_decap_8 FILLER_27_931 ();
 sg13g2_decap_8 FILLER_27_938 ();
 sg13g2_decap_8 FILLER_27_945 ();
 sg13g2_decap_8 FILLER_27_952 ();
 sg13g2_decap_8 FILLER_27_959 ();
 sg13g2_decap_8 FILLER_27_966 ();
 sg13g2_decap_8 FILLER_27_973 ();
 sg13g2_decap_8 FILLER_27_980 ();
 sg13g2_decap_8 FILLER_27_987 ();
 sg13g2_decap_8 FILLER_27_994 ();
 sg13g2_decap_8 FILLER_27_1001 ();
 sg13g2_decap_8 FILLER_27_1008 ();
 sg13g2_decap_8 FILLER_27_1015 ();
 sg13g2_decap_8 FILLER_27_1022 ();
 sg13g2_decap_8 FILLER_28_4 ();
 sg13g2_decap_8 FILLER_28_11 ();
 sg13g2_decap_8 FILLER_28_18 ();
 sg13g2_decap_8 FILLER_28_25 ();
 sg13g2_decap_8 FILLER_28_32 ();
 sg13g2_decap_8 FILLER_28_39 ();
 sg13g2_decap_8 FILLER_28_46 ();
 sg13g2_decap_8 FILLER_28_53 ();
 sg13g2_decap_8 FILLER_28_60 ();
 sg13g2_decap_8 FILLER_28_67 ();
 sg13g2_decap_8 FILLER_28_74 ();
 sg13g2_decap_8 FILLER_28_81 ();
 sg13g2_decap_8 FILLER_28_88 ();
 sg13g2_decap_8 FILLER_28_95 ();
 sg13g2_decap_8 FILLER_28_102 ();
 sg13g2_decap_8 FILLER_28_109 ();
 sg13g2_decap_8 FILLER_28_116 ();
 sg13g2_decap_8 FILLER_28_123 ();
 sg13g2_decap_8 FILLER_28_130 ();
 sg13g2_decap_8 FILLER_28_137 ();
 sg13g2_decap_4 FILLER_28_144 ();
 sg13g2_fill_1 FILLER_28_148 ();
 sg13g2_decap_8 FILLER_28_176 ();
 sg13g2_decap_8 FILLER_28_183 ();
 sg13g2_decap_8 FILLER_28_190 ();
 sg13g2_decap_8 FILLER_28_197 ();
 sg13g2_decap_8 FILLER_28_204 ();
 sg13g2_decap_8 FILLER_28_211 ();
 sg13g2_decap_8 FILLER_28_218 ();
 sg13g2_decap_8 FILLER_28_225 ();
 sg13g2_decap_8 FILLER_28_232 ();
 sg13g2_decap_4 FILLER_28_239 ();
 sg13g2_fill_2 FILLER_28_243 ();
 sg13g2_decap_8 FILLER_28_272 ();
 sg13g2_decap_8 FILLER_28_279 ();
 sg13g2_decap_4 FILLER_28_286 ();
 sg13g2_fill_2 FILLER_28_290 ();
 sg13g2_decap_8 FILLER_28_300 ();
 sg13g2_decap_8 FILLER_28_307 ();
 sg13g2_decap_8 FILLER_28_314 ();
 sg13g2_decap_8 FILLER_28_321 ();
 sg13g2_fill_2 FILLER_28_328 ();
 sg13g2_fill_1 FILLER_28_330 ();
 sg13g2_decap_8 FILLER_28_335 ();
 sg13g2_decap_4 FILLER_28_342 ();
 sg13g2_fill_2 FILLER_28_346 ();
 sg13g2_decap_8 FILLER_28_368 ();
 sg13g2_decap_8 FILLER_28_375 ();
 sg13g2_decap_8 FILLER_28_382 ();
 sg13g2_decap_8 FILLER_28_389 ();
 sg13g2_decap_4 FILLER_28_396 ();
 sg13g2_fill_1 FILLER_28_400 ();
 sg13g2_decap_8 FILLER_28_428 ();
 sg13g2_decap_8 FILLER_28_435 ();
 sg13g2_decap_8 FILLER_28_442 ();
 sg13g2_decap_8 FILLER_28_449 ();
 sg13g2_decap_8 FILLER_28_456 ();
 sg13g2_decap_8 FILLER_28_463 ();
 sg13g2_decap_8 FILLER_28_470 ();
 sg13g2_decap_8 FILLER_28_477 ();
 sg13g2_decap_8 FILLER_28_484 ();
 sg13g2_decap_8 FILLER_28_491 ();
 sg13g2_decap_8 FILLER_28_498 ();
 sg13g2_decap_8 FILLER_28_505 ();
 sg13g2_decap_8 FILLER_28_512 ();
 sg13g2_decap_8 FILLER_28_519 ();
 sg13g2_decap_8 FILLER_28_526 ();
 sg13g2_decap_8 FILLER_28_533 ();
 sg13g2_decap_8 FILLER_28_540 ();
 sg13g2_decap_8 FILLER_28_547 ();
 sg13g2_decap_8 FILLER_28_554 ();
 sg13g2_decap_8 FILLER_28_561 ();
 sg13g2_decap_8 FILLER_28_568 ();
 sg13g2_decap_8 FILLER_28_575 ();
 sg13g2_decap_8 FILLER_28_582 ();
 sg13g2_decap_8 FILLER_28_589 ();
 sg13g2_decap_8 FILLER_28_596 ();
 sg13g2_decap_8 FILLER_28_603 ();
 sg13g2_decap_8 FILLER_28_610 ();
 sg13g2_decap_8 FILLER_28_617 ();
 sg13g2_decap_8 FILLER_28_624 ();
 sg13g2_decap_8 FILLER_28_631 ();
 sg13g2_decap_8 FILLER_28_638 ();
 sg13g2_decap_8 FILLER_28_645 ();
 sg13g2_decap_8 FILLER_28_652 ();
 sg13g2_decap_8 FILLER_28_659 ();
 sg13g2_decap_8 FILLER_28_666 ();
 sg13g2_decap_8 FILLER_28_673 ();
 sg13g2_decap_8 FILLER_28_680 ();
 sg13g2_decap_8 FILLER_28_687 ();
 sg13g2_decap_8 FILLER_28_694 ();
 sg13g2_decap_8 FILLER_28_701 ();
 sg13g2_decap_8 FILLER_28_708 ();
 sg13g2_decap_8 FILLER_28_715 ();
 sg13g2_decap_8 FILLER_28_722 ();
 sg13g2_decap_8 FILLER_28_729 ();
 sg13g2_decap_8 FILLER_28_736 ();
 sg13g2_decap_8 FILLER_28_743 ();
 sg13g2_decap_8 FILLER_28_750 ();
 sg13g2_decap_8 FILLER_28_757 ();
 sg13g2_decap_8 FILLER_28_764 ();
 sg13g2_decap_8 FILLER_28_771 ();
 sg13g2_decap_8 FILLER_28_778 ();
 sg13g2_decap_8 FILLER_28_785 ();
 sg13g2_decap_8 FILLER_28_792 ();
 sg13g2_decap_8 FILLER_28_799 ();
 sg13g2_decap_8 FILLER_28_806 ();
 sg13g2_decap_8 FILLER_28_813 ();
 sg13g2_decap_8 FILLER_28_820 ();
 sg13g2_decap_8 FILLER_28_827 ();
 sg13g2_decap_8 FILLER_28_834 ();
 sg13g2_decap_8 FILLER_28_841 ();
 sg13g2_decap_8 FILLER_28_848 ();
 sg13g2_decap_8 FILLER_28_855 ();
 sg13g2_decap_8 FILLER_28_862 ();
 sg13g2_decap_8 FILLER_28_869 ();
 sg13g2_decap_8 FILLER_28_876 ();
 sg13g2_decap_8 FILLER_28_883 ();
 sg13g2_decap_8 FILLER_28_890 ();
 sg13g2_decap_8 FILLER_28_897 ();
 sg13g2_decap_8 FILLER_28_904 ();
 sg13g2_decap_8 FILLER_28_911 ();
 sg13g2_decap_8 FILLER_28_918 ();
 sg13g2_decap_8 FILLER_28_925 ();
 sg13g2_decap_8 FILLER_28_932 ();
 sg13g2_decap_8 FILLER_28_939 ();
 sg13g2_decap_8 FILLER_28_946 ();
 sg13g2_decap_8 FILLER_28_953 ();
 sg13g2_decap_8 FILLER_28_960 ();
 sg13g2_decap_8 FILLER_28_967 ();
 sg13g2_decap_8 FILLER_28_974 ();
 sg13g2_decap_8 FILLER_28_981 ();
 sg13g2_decap_8 FILLER_28_988 ();
 sg13g2_decap_8 FILLER_28_995 ();
 sg13g2_decap_8 FILLER_28_1002 ();
 sg13g2_decap_8 FILLER_28_1009 ();
 sg13g2_decap_8 FILLER_28_1016 ();
 sg13g2_decap_4 FILLER_28_1023 ();
 sg13g2_fill_2 FILLER_28_1027 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_decap_8 FILLER_29_105 ();
 sg13g2_decap_8 FILLER_29_112 ();
 sg13g2_decap_8 FILLER_29_119 ();
 sg13g2_decap_8 FILLER_29_126 ();
 sg13g2_decap_8 FILLER_29_133 ();
 sg13g2_decap_8 FILLER_29_140 ();
 sg13g2_decap_8 FILLER_29_147 ();
 sg13g2_decap_8 FILLER_29_154 ();
 sg13g2_decap_8 FILLER_29_161 ();
 sg13g2_decap_8 FILLER_29_168 ();
 sg13g2_decap_8 FILLER_29_175 ();
 sg13g2_decap_8 FILLER_29_182 ();
 sg13g2_decap_4 FILLER_29_189 ();
 sg13g2_fill_2 FILLER_29_193 ();
 sg13g2_decap_8 FILLER_29_222 ();
 sg13g2_decap_8 FILLER_29_229 ();
 sg13g2_decap_8 FILLER_29_236 ();
 sg13g2_decap_8 FILLER_29_243 ();
 sg13g2_decap_8 FILLER_29_250 ();
 sg13g2_decap_8 FILLER_29_257 ();
 sg13g2_decap_8 FILLER_29_264 ();
 sg13g2_decap_8 FILLER_29_271 ();
 sg13g2_decap_8 FILLER_29_278 ();
 sg13g2_decap_4 FILLER_29_285 ();
 sg13g2_fill_2 FILLER_29_289 ();
 sg13g2_decap_8 FILLER_29_296 ();
 sg13g2_decap_8 FILLER_29_303 ();
 sg13g2_decap_8 FILLER_29_310 ();
 sg13g2_decap_8 FILLER_29_317 ();
 sg13g2_decap_8 FILLER_29_324 ();
 sg13g2_decap_8 FILLER_29_331 ();
 sg13g2_decap_8 FILLER_29_338 ();
 sg13g2_fill_2 FILLER_29_345 ();
 sg13g2_fill_1 FILLER_29_347 ();
 sg13g2_decap_8 FILLER_29_375 ();
 sg13g2_decap_8 FILLER_29_382 ();
 sg13g2_decap_8 FILLER_29_389 ();
 sg13g2_decap_8 FILLER_29_396 ();
 sg13g2_decap_8 FILLER_29_403 ();
 sg13g2_decap_8 FILLER_29_410 ();
 sg13g2_decap_8 FILLER_29_417 ();
 sg13g2_decap_8 FILLER_29_424 ();
 sg13g2_decap_8 FILLER_29_431 ();
 sg13g2_decap_8 FILLER_29_438 ();
 sg13g2_decap_8 FILLER_29_445 ();
 sg13g2_decap_8 FILLER_29_452 ();
 sg13g2_decap_8 FILLER_29_459 ();
 sg13g2_decap_8 FILLER_29_466 ();
 sg13g2_decap_8 FILLER_29_473 ();
 sg13g2_decap_8 FILLER_29_480 ();
 sg13g2_decap_8 FILLER_29_487 ();
 sg13g2_decap_8 FILLER_29_494 ();
 sg13g2_decap_8 FILLER_29_501 ();
 sg13g2_decap_8 FILLER_29_508 ();
 sg13g2_decap_8 FILLER_29_515 ();
 sg13g2_decap_8 FILLER_29_522 ();
 sg13g2_decap_8 FILLER_29_529 ();
 sg13g2_decap_8 FILLER_29_536 ();
 sg13g2_decap_8 FILLER_29_543 ();
 sg13g2_decap_8 FILLER_29_550 ();
 sg13g2_decap_8 FILLER_29_557 ();
 sg13g2_decap_8 FILLER_29_564 ();
 sg13g2_decap_8 FILLER_29_571 ();
 sg13g2_decap_8 FILLER_29_578 ();
 sg13g2_decap_8 FILLER_29_585 ();
 sg13g2_decap_8 FILLER_29_592 ();
 sg13g2_decap_8 FILLER_29_599 ();
 sg13g2_decap_8 FILLER_29_606 ();
 sg13g2_decap_8 FILLER_29_613 ();
 sg13g2_decap_8 FILLER_29_620 ();
 sg13g2_decap_8 FILLER_29_627 ();
 sg13g2_decap_8 FILLER_29_634 ();
 sg13g2_decap_8 FILLER_29_641 ();
 sg13g2_decap_8 FILLER_29_648 ();
 sg13g2_decap_8 FILLER_29_655 ();
 sg13g2_decap_8 FILLER_29_662 ();
 sg13g2_decap_8 FILLER_29_669 ();
 sg13g2_decap_8 FILLER_29_676 ();
 sg13g2_decap_8 FILLER_29_683 ();
 sg13g2_decap_8 FILLER_29_690 ();
 sg13g2_decap_8 FILLER_29_697 ();
 sg13g2_decap_8 FILLER_29_704 ();
 sg13g2_decap_8 FILLER_29_711 ();
 sg13g2_decap_8 FILLER_29_718 ();
 sg13g2_decap_8 FILLER_29_725 ();
 sg13g2_decap_8 FILLER_29_732 ();
 sg13g2_decap_8 FILLER_29_739 ();
 sg13g2_decap_8 FILLER_29_746 ();
 sg13g2_decap_8 FILLER_29_753 ();
 sg13g2_decap_8 FILLER_29_760 ();
 sg13g2_decap_8 FILLER_29_767 ();
 sg13g2_decap_8 FILLER_29_774 ();
 sg13g2_decap_8 FILLER_29_781 ();
 sg13g2_decap_8 FILLER_29_788 ();
 sg13g2_decap_8 FILLER_29_795 ();
 sg13g2_decap_8 FILLER_29_802 ();
 sg13g2_decap_8 FILLER_29_809 ();
 sg13g2_decap_8 FILLER_29_816 ();
 sg13g2_decap_8 FILLER_29_823 ();
 sg13g2_decap_8 FILLER_29_830 ();
 sg13g2_decap_8 FILLER_29_837 ();
 sg13g2_decap_8 FILLER_29_844 ();
 sg13g2_decap_8 FILLER_29_851 ();
 sg13g2_decap_8 FILLER_29_858 ();
 sg13g2_decap_8 FILLER_29_865 ();
 sg13g2_decap_8 FILLER_29_872 ();
 sg13g2_decap_8 FILLER_29_879 ();
 sg13g2_decap_8 FILLER_29_886 ();
 sg13g2_decap_8 FILLER_29_893 ();
 sg13g2_decap_8 FILLER_29_900 ();
 sg13g2_decap_8 FILLER_29_907 ();
 sg13g2_decap_8 FILLER_29_914 ();
 sg13g2_decap_8 FILLER_29_921 ();
 sg13g2_decap_8 FILLER_29_928 ();
 sg13g2_decap_8 FILLER_29_935 ();
 sg13g2_decap_8 FILLER_29_942 ();
 sg13g2_decap_8 FILLER_29_949 ();
 sg13g2_decap_8 FILLER_29_956 ();
 sg13g2_decap_8 FILLER_29_963 ();
 sg13g2_decap_8 FILLER_29_970 ();
 sg13g2_decap_8 FILLER_29_977 ();
 sg13g2_decap_8 FILLER_29_984 ();
 sg13g2_decap_8 FILLER_29_991 ();
 sg13g2_decap_8 FILLER_29_998 ();
 sg13g2_decap_8 FILLER_29_1005 ();
 sg13g2_decap_8 FILLER_29_1012 ();
 sg13g2_decap_8 FILLER_29_1019 ();
 sg13g2_fill_2 FILLER_29_1026 ();
 sg13g2_fill_1 FILLER_29_1028 ();
 sg13g2_decap_8 FILLER_30_5 ();
 sg13g2_decap_8 FILLER_30_12 ();
 sg13g2_decap_8 FILLER_30_19 ();
 sg13g2_decap_8 FILLER_30_26 ();
 sg13g2_decap_8 FILLER_30_33 ();
 sg13g2_decap_8 FILLER_30_40 ();
 sg13g2_decap_8 FILLER_30_47 ();
 sg13g2_decap_8 FILLER_30_54 ();
 sg13g2_decap_8 FILLER_30_61 ();
 sg13g2_decap_8 FILLER_30_68 ();
 sg13g2_decap_8 FILLER_30_75 ();
 sg13g2_decap_8 FILLER_30_82 ();
 sg13g2_decap_8 FILLER_30_89 ();
 sg13g2_decap_8 FILLER_30_96 ();
 sg13g2_decap_8 FILLER_30_103 ();
 sg13g2_decap_8 FILLER_30_110 ();
 sg13g2_decap_8 FILLER_30_117 ();
 sg13g2_decap_8 FILLER_30_124 ();
 sg13g2_decap_8 FILLER_30_131 ();
 sg13g2_decap_8 FILLER_30_138 ();
 sg13g2_decap_8 FILLER_30_145 ();
 sg13g2_decap_8 FILLER_30_152 ();
 sg13g2_decap_8 FILLER_30_159 ();
 sg13g2_decap_8 FILLER_30_166 ();
 sg13g2_decap_8 FILLER_30_173 ();
 sg13g2_decap_8 FILLER_30_180 ();
 sg13g2_decap_8 FILLER_30_187 ();
 sg13g2_decap_8 FILLER_30_194 ();
 sg13g2_decap_8 FILLER_30_201 ();
 sg13g2_decap_8 FILLER_30_208 ();
 sg13g2_decap_8 FILLER_30_215 ();
 sg13g2_decap_8 FILLER_30_222 ();
 sg13g2_decap_8 FILLER_30_229 ();
 sg13g2_decap_8 FILLER_30_236 ();
 sg13g2_decap_8 FILLER_30_243 ();
 sg13g2_decap_8 FILLER_30_250 ();
 sg13g2_decap_8 FILLER_30_257 ();
 sg13g2_decap_8 FILLER_30_264 ();
 sg13g2_decap_8 FILLER_30_271 ();
 sg13g2_decap_8 FILLER_30_278 ();
 sg13g2_decap_8 FILLER_30_285 ();
 sg13g2_fill_2 FILLER_30_292 ();
 sg13g2_decap_8 FILLER_30_297 ();
 sg13g2_decap_8 FILLER_30_304 ();
 sg13g2_decap_8 FILLER_30_311 ();
 sg13g2_decap_8 FILLER_30_318 ();
 sg13g2_decap_8 FILLER_30_325 ();
 sg13g2_fill_2 FILLER_30_332 ();
 sg13g2_fill_1 FILLER_30_334 ();
 sg13g2_decap_8 FILLER_30_352 ();
 sg13g2_decap_8 FILLER_30_359 ();
 sg13g2_decap_8 FILLER_30_366 ();
 sg13g2_decap_8 FILLER_30_373 ();
 sg13g2_decap_8 FILLER_30_380 ();
 sg13g2_decap_8 FILLER_30_387 ();
 sg13g2_decap_8 FILLER_30_394 ();
 sg13g2_decap_8 FILLER_30_401 ();
 sg13g2_decap_8 FILLER_30_408 ();
 sg13g2_decap_8 FILLER_30_415 ();
 sg13g2_decap_8 FILLER_30_422 ();
 sg13g2_decap_8 FILLER_30_429 ();
 sg13g2_decap_8 FILLER_30_436 ();
 sg13g2_decap_8 FILLER_30_443 ();
 sg13g2_decap_8 FILLER_30_450 ();
 sg13g2_decap_8 FILLER_30_457 ();
 sg13g2_decap_8 FILLER_30_464 ();
 sg13g2_decap_8 FILLER_30_471 ();
 sg13g2_decap_8 FILLER_30_478 ();
 sg13g2_decap_8 FILLER_30_485 ();
 sg13g2_decap_8 FILLER_30_492 ();
 sg13g2_decap_8 FILLER_30_499 ();
 sg13g2_decap_8 FILLER_30_506 ();
 sg13g2_decap_8 FILLER_30_513 ();
 sg13g2_decap_8 FILLER_30_520 ();
 sg13g2_decap_8 FILLER_30_527 ();
 sg13g2_decap_8 FILLER_30_534 ();
 sg13g2_decap_8 FILLER_30_541 ();
 sg13g2_decap_8 FILLER_30_548 ();
 sg13g2_decap_8 FILLER_30_555 ();
 sg13g2_decap_8 FILLER_30_562 ();
 sg13g2_decap_8 FILLER_30_569 ();
 sg13g2_decap_8 FILLER_30_576 ();
 sg13g2_decap_8 FILLER_30_583 ();
 sg13g2_decap_8 FILLER_30_590 ();
 sg13g2_decap_8 FILLER_30_597 ();
 sg13g2_decap_8 FILLER_30_604 ();
 sg13g2_decap_8 FILLER_30_611 ();
 sg13g2_decap_8 FILLER_30_618 ();
 sg13g2_decap_8 FILLER_30_625 ();
 sg13g2_decap_8 FILLER_30_632 ();
 sg13g2_decap_8 FILLER_30_639 ();
 sg13g2_decap_8 FILLER_30_646 ();
 sg13g2_decap_8 FILLER_30_653 ();
 sg13g2_decap_8 FILLER_30_660 ();
 sg13g2_decap_8 FILLER_30_667 ();
 sg13g2_decap_8 FILLER_30_674 ();
 sg13g2_decap_8 FILLER_30_681 ();
 sg13g2_decap_8 FILLER_30_688 ();
 sg13g2_decap_8 FILLER_30_695 ();
 sg13g2_decap_8 FILLER_30_702 ();
 sg13g2_decap_8 FILLER_30_709 ();
 sg13g2_decap_8 FILLER_30_716 ();
 sg13g2_decap_8 FILLER_30_723 ();
 sg13g2_decap_8 FILLER_30_730 ();
 sg13g2_decap_8 FILLER_30_737 ();
 sg13g2_decap_8 FILLER_30_744 ();
 sg13g2_decap_8 FILLER_30_751 ();
 sg13g2_decap_8 FILLER_30_758 ();
 sg13g2_decap_8 FILLER_30_765 ();
 sg13g2_decap_8 FILLER_30_772 ();
 sg13g2_decap_8 FILLER_30_779 ();
 sg13g2_decap_8 FILLER_30_786 ();
 sg13g2_decap_8 FILLER_30_793 ();
 sg13g2_decap_8 FILLER_30_800 ();
 sg13g2_decap_8 FILLER_30_807 ();
 sg13g2_decap_8 FILLER_30_814 ();
 sg13g2_decap_8 FILLER_30_821 ();
 sg13g2_decap_8 FILLER_30_828 ();
 sg13g2_decap_8 FILLER_30_835 ();
 sg13g2_decap_8 FILLER_30_842 ();
 sg13g2_decap_8 FILLER_30_849 ();
 sg13g2_decap_8 FILLER_30_856 ();
 sg13g2_decap_8 FILLER_30_863 ();
 sg13g2_decap_8 FILLER_30_870 ();
 sg13g2_decap_8 FILLER_30_877 ();
 sg13g2_decap_8 FILLER_30_884 ();
 sg13g2_decap_8 FILLER_30_891 ();
 sg13g2_decap_8 FILLER_30_898 ();
 sg13g2_decap_8 FILLER_30_905 ();
 sg13g2_decap_8 FILLER_30_912 ();
 sg13g2_decap_8 FILLER_30_919 ();
 sg13g2_decap_8 FILLER_30_926 ();
 sg13g2_decap_8 FILLER_30_933 ();
 sg13g2_decap_8 FILLER_30_940 ();
 sg13g2_decap_8 FILLER_30_947 ();
 sg13g2_decap_8 FILLER_30_954 ();
 sg13g2_decap_8 FILLER_30_961 ();
 sg13g2_decap_8 FILLER_30_968 ();
 sg13g2_decap_8 FILLER_30_975 ();
 sg13g2_decap_8 FILLER_30_982 ();
 sg13g2_decap_8 FILLER_30_989 ();
 sg13g2_decap_8 FILLER_30_996 ();
 sg13g2_decap_8 FILLER_30_1003 ();
 sg13g2_decap_8 FILLER_30_1010 ();
 sg13g2_decap_8 FILLER_30_1017 ();
 sg13g2_decap_4 FILLER_30_1024 ();
 sg13g2_fill_1 FILLER_30_1028 ();
 sg13g2_decap_8 FILLER_31_5 ();
 sg13g2_decap_8 FILLER_31_12 ();
 sg13g2_decap_8 FILLER_31_19 ();
 sg13g2_decap_8 FILLER_31_26 ();
 sg13g2_decap_8 FILLER_31_33 ();
 sg13g2_decap_8 FILLER_31_40 ();
 sg13g2_decap_8 FILLER_31_47 ();
 sg13g2_decap_8 FILLER_31_54 ();
 sg13g2_decap_8 FILLER_31_61 ();
 sg13g2_decap_8 FILLER_31_68 ();
 sg13g2_decap_8 FILLER_31_75 ();
 sg13g2_decap_8 FILLER_31_82 ();
 sg13g2_decap_8 FILLER_31_89 ();
 sg13g2_decap_8 FILLER_31_96 ();
 sg13g2_decap_8 FILLER_31_103 ();
 sg13g2_decap_8 FILLER_31_110 ();
 sg13g2_decap_8 FILLER_31_117 ();
 sg13g2_decap_8 FILLER_31_124 ();
 sg13g2_decap_8 FILLER_31_131 ();
 sg13g2_decap_8 FILLER_31_138 ();
 sg13g2_decap_8 FILLER_31_145 ();
 sg13g2_decap_8 FILLER_31_152 ();
 sg13g2_decap_8 FILLER_31_159 ();
 sg13g2_decap_8 FILLER_31_166 ();
 sg13g2_decap_8 FILLER_31_173 ();
 sg13g2_decap_8 FILLER_31_180 ();
 sg13g2_decap_8 FILLER_31_187 ();
 sg13g2_decap_8 FILLER_31_194 ();
 sg13g2_decap_8 FILLER_31_201 ();
 sg13g2_decap_8 FILLER_31_208 ();
 sg13g2_decap_8 FILLER_31_215 ();
 sg13g2_decap_8 FILLER_31_222 ();
 sg13g2_decap_8 FILLER_31_246 ();
 sg13g2_decap_8 FILLER_31_253 ();
 sg13g2_decap_8 FILLER_31_260 ();
 sg13g2_decap_8 FILLER_31_267 ();
 sg13g2_decap_8 FILLER_31_274 ();
 sg13g2_decap_8 FILLER_31_281 ();
 sg13g2_decap_8 FILLER_31_288 ();
 sg13g2_decap_8 FILLER_31_295 ();
 sg13g2_decap_8 FILLER_31_309 ();
 sg13g2_decap_8 FILLER_31_316 ();
 sg13g2_decap_8 FILLER_31_323 ();
 sg13g2_decap_8 FILLER_31_330 ();
 sg13g2_decap_8 FILLER_31_337 ();
 sg13g2_decap_8 FILLER_31_344 ();
 sg13g2_decap_8 FILLER_31_351 ();
 sg13g2_decap_8 FILLER_31_358 ();
 sg13g2_decap_8 FILLER_31_365 ();
 sg13g2_decap_8 FILLER_31_372 ();
 sg13g2_decap_8 FILLER_31_379 ();
 sg13g2_decap_8 FILLER_31_386 ();
 sg13g2_decap_8 FILLER_31_393 ();
 sg13g2_decap_8 FILLER_31_400 ();
 sg13g2_decap_8 FILLER_31_407 ();
 sg13g2_decap_8 FILLER_31_414 ();
 sg13g2_decap_8 FILLER_31_421 ();
 sg13g2_decap_8 FILLER_31_428 ();
 sg13g2_decap_8 FILLER_31_435 ();
 sg13g2_decap_8 FILLER_31_442 ();
 sg13g2_decap_8 FILLER_31_449 ();
 sg13g2_decap_8 FILLER_31_456 ();
 sg13g2_decap_8 FILLER_31_463 ();
 sg13g2_decap_8 FILLER_31_470 ();
 sg13g2_decap_8 FILLER_31_477 ();
 sg13g2_decap_8 FILLER_31_484 ();
 sg13g2_decap_8 FILLER_31_491 ();
 sg13g2_decap_8 FILLER_31_498 ();
 sg13g2_decap_8 FILLER_31_505 ();
 sg13g2_decap_8 FILLER_31_512 ();
 sg13g2_decap_8 FILLER_31_519 ();
 sg13g2_decap_8 FILLER_31_526 ();
 sg13g2_decap_8 FILLER_31_533 ();
 sg13g2_decap_8 FILLER_31_540 ();
 sg13g2_decap_8 FILLER_31_547 ();
 sg13g2_decap_8 FILLER_31_554 ();
 sg13g2_decap_8 FILLER_31_561 ();
 sg13g2_decap_8 FILLER_31_568 ();
 sg13g2_decap_8 FILLER_31_575 ();
 sg13g2_decap_8 FILLER_31_582 ();
 sg13g2_decap_8 FILLER_31_589 ();
 sg13g2_decap_8 FILLER_31_596 ();
 sg13g2_decap_8 FILLER_31_603 ();
 sg13g2_decap_8 FILLER_31_610 ();
 sg13g2_decap_8 FILLER_31_617 ();
 sg13g2_decap_8 FILLER_31_624 ();
 sg13g2_decap_8 FILLER_31_631 ();
 sg13g2_decap_8 FILLER_31_638 ();
 sg13g2_decap_8 FILLER_31_645 ();
 sg13g2_decap_8 FILLER_31_652 ();
 sg13g2_decap_8 FILLER_31_659 ();
 sg13g2_decap_8 FILLER_31_666 ();
 sg13g2_decap_8 FILLER_31_673 ();
 sg13g2_decap_8 FILLER_31_680 ();
 sg13g2_decap_8 FILLER_31_687 ();
 sg13g2_decap_8 FILLER_31_694 ();
 sg13g2_decap_8 FILLER_31_701 ();
 sg13g2_decap_8 FILLER_31_708 ();
 sg13g2_decap_8 FILLER_31_715 ();
 sg13g2_decap_8 FILLER_31_722 ();
 sg13g2_decap_8 FILLER_31_729 ();
 sg13g2_decap_8 FILLER_31_736 ();
 sg13g2_decap_8 FILLER_31_743 ();
 sg13g2_decap_8 FILLER_31_750 ();
 sg13g2_decap_8 FILLER_31_757 ();
 sg13g2_decap_8 FILLER_31_764 ();
 sg13g2_decap_8 FILLER_31_771 ();
 sg13g2_decap_8 FILLER_31_778 ();
 sg13g2_decap_8 FILLER_31_785 ();
 sg13g2_decap_8 FILLER_31_792 ();
 sg13g2_decap_8 FILLER_31_799 ();
 sg13g2_decap_8 FILLER_31_806 ();
 sg13g2_decap_8 FILLER_31_813 ();
 sg13g2_decap_8 FILLER_31_820 ();
 sg13g2_decap_8 FILLER_31_827 ();
 sg13g2_decap_8 FILLER_31_834 ();
 sg13g2_decap_8 FILLER_31_841 ();
 sg13g2_decap_8 FILLER_31_848 ();
 sg13g2_decap_8 FILLER_31_855 ();
 sg13g2_decap_8 FILLER_31_862 ();
 sg13g2_decap_8 FILLER_31_869 ();
 sg13g2_decap_8 FILLER_31_876 ();
 sg13g2_decap_8 FILLER_31_883 ();
 sg13g2_decap_8 FILLER_31_890 ();
 sg13g2_decap_8 FILLER_31_897 ();
 sg13g2_decap_8 FILLER_31_904 ();
 sg13g2_decap_8 FILLER_31_911 ();
 sg13g2_decap_8 FILLER_31_918 ();
 sg13g2_decap_8 FILLER_31_925 ();
 sg13g2_decap_8 FILLER_31_932 ();
 sg13g2_decap_8 FILLER_31_939 ();
 sg13g2_decap_8 FILLER_31_946 ();
 sg13g2_decap_8 FILLER_31_953 ();
 sg13g2_decap_8 FILLER_31_960 ();
 sg13g2_decap_8 FILLER_31_967 ();
 sg13g2_decap_8 FILLER_31_974 ();
 sg13g2_decap_8 FILLER_31_981 ();
 sg13g2_decap_8 FILLER_31_988 ();
 sg13g2_decap_8 FILLER_31_995 ();
 sg13g2_decap_8 FILLER_31_1002 ();
 sg13g2_decap_8 FILLER_31_1009 ();
 sg13g2_decap_8 FILLER_31_1016 ();
 sg13g2_decap_4 FILLER_31_1023 ();
 sg13g2_fill_2 FILLER_31_1027 ();
 sg13g2_decap_8 FILLER_32_5 ();
 sg13g2_decap_8 FILLER_32_12 ();
 sg13g2_decap_8 FILLER_32_19 ();
 sg13g2_decap_8 FILLER_32_26 ();
 sg13g2_decap_8 FILLER_32_33 ();
 sg13g2_decap_8 FILLER_32_40 ();
 sg13g2_decap_8 FILLER_32_47 ();
 sg13g2_decap_8 FILLER_32_54 ();
 sg13g2_decap_8 FILLER_32_61 ();
 sg13g2_decap_8 FILLER_32_68 ();
 sg13g2_decap_8 FILLER_32_75 ();
 sg13g2_decap_8 FILLER_32_82 ();
 sg13g2_decap_8 FILLER_32_89 ();
 sg13g2_decap_8 FILLER_32_96 ();
 sg13g2_decap_8 FILLER_32_103 ();
 sg13g2_decap_8 FILLER_32_110 ();
 sg13g2_decap_8 FILLER_32_117 ();
 sg13g2_decap_8 FILLER_32_124 ();
 sg13g2_decap_8 FILLER_32_131 ();
 sg13g2_decap_8 FILLER_32_138 ();
 sg13g2_decap_8 FILLER_32_145 ();
 sg13g2_decap_8 FILLER_32_152 ();
 sg13g2_decap_8 FILLER_32_159 ();
 sg13g2_decap_8 FILLER_32_166 ();
 sg13g2_decap_8 FILLER_32_173 ();
 sg13g2_decap_8 FILLER_32_180 ();
 sg13g2_decap_8 FILLER_32_187 ();
 sg13g2_decap_8 FILLER_32_194 ();
 sg13g2_decap_8 FILLER_32_201 ();
 sg13g2_decap_8 FILLER_32_208 ();
 sg13g2_decap_8 FILLER_32_215 ();
 sg13g2_decap_8 FILLER_32_222 ();
 sg13g2_decap_8 FILLER_32_229 ();
 sg13g2_decap_8 FILLER_32_236 ();
 sg13g2_decap_8 FILLER_32_243 ();
 sg13g2_decap_8 FILLER_32_250 ();
 sg13g2_decap_8 FILLER_32_257 ();
 sg13g2_decap_8 FILLER_32_264 ();
 sg13g2_decap_8 FILLER_32_271 ();
 sg13g2_decap_8 FILLER_32_278 ();
 sg13g2_fill_2 FILLER_32_285 ();
 sg13g2_decap_8 FILLER_32_292 ();
 sg13g2_decap_8 FILLER_32_299 ();
 sg13g2_decap_8 FILLER_32_306 ();
 sg13g2_decap_8 FILLER_32_313 ();
 sg13g2_decap_8 FILLER_32_320 ();
 sg13g2_decap_8 FILLER_32_327 ();
 sg13g2_decap_8 FILLER_32_334 ();
 sg13g2_decap_8 FILLER_32_341 ();
 sg13g2_decap_8 FILLER_32_348 ();
 sg13g2_decap_8 FILLER_32_355 ();
 sg13g2_decap_8 FILLER_32_362 ();
 sg13g2_decap_8 FILLER_32_369 ();
 sg13g2_decap_8 FILLER_32_376 ();
 sg13g2_decap_8 FILLER_32_383 ();
 sg13g2_decap_8 FILLER_32_390 ();
 sg13g2_decap_8 FILLER_32_397 ();
 sg13g2_decap_8 FILLER_32_404 ();
 sg13g2_decap_8 FILLER_32_411 ();
 sg13g2_decap_8 FILLER_32_418 ();
 sg13g2_decap_8 FILLER_32_425 ();
 sg13g2_decap_8 FILLER_32_432 ();
 sg13g2_decap_8 FILLER_32_439 ();
 sg13g2_decap_8 FILLER_32_446 ();
 sg13g2_decap_8 FILLER_32_453 ();
 sg13g2_decap_8 FILLER_32_460 ();
 sg13g2_decap_8 FILLER_32_467 ();
 sg13g2_decap_8 FILLER_32_474 ();
 sg13g2_decap_8 FILLER_32_481 ();
 sg13g2_decap_8 FILLER_32_488 ();
 sg13g2_decap_8 FILLER_32_495 ();
 sg13g2_decap_8 FILLER_32_502 ();
 sg13g2_decap_8 FILLER_32_509 ();
 sg13g2_decap_8 FILLER_32_516 ();
 sg13g2_decap_8 FILLER_32_523 ();
 sg13g2_decap_8 FILLER_32_530 ();
 sg13g2_decap_8 FILLER_32_537 ();
 sg13g2_decap_8 FILLER_32_544 ();
 sg13g2_decap_8 FILLER_32_551 ();
 sg13g2_decap_8 FILLER_32_558 ();
 sg13g2_decap_8 FILLER_32_565 ();
 sg13g2_decap_8 FILLER_32_572 ();
 sg13g2_decap_8 FILLER_32_579 ();
 sg13g2_decap_8 FILLER_32_586 ();
 sg13g2_decap_8 FILLER_32_593 ();
 sg13g2_decap_8 FILLER_32_600 ();
 sg13g2_decap_8 FILLER_32_607 ();
 sg13g2_decap_8 FILLER_32_614 ();
 sg13g2_decap_8 FILLER_32_621 ();
 sg13g2_decap_8 FILLER_32_628 ();
 sg13g2_decap_8 FILLER_32_635 ();
 sg13g2_decap_8 FILLER_32_642 ();
 sg13g2_decap_8 FILLER_32_649 ();
 sg13g2_decap_8 FILLER_32_656 ();
 sg13g2_decap_8 FILLER_32_663 ();
 sg13g2_decap_8 FILLER_32_670 ();
 sg13g2_decap_8 FILLER_32_677 ();
 sg13g2_decap_8 FILLER_32_684 ();
 sg13g2_decap_8 FILLER_32_691 ();
 sg13g2_decap_8 FILLER_32_698 ();
 sg13g2_decap_8 FILLER_32_705 ();
 sg13g2_decap_8 FILLER_32_712 ();
 sg13g2_decap_8 FILLER_32_719 ();
 sg13g2_decap_8 FILLER_32_726 ();
 sg13g2_decap_8 FILLER_32_733 ();
 sg13g2_decap_8 FILLER_32_740 ();
 sg13g2_decap_8 FILLER_32_747 ();
 sg13g2_decap_8 FILLER_32_754 ();
 sg13g2_decap_8 FILLER_32_761 ();
 sg13g2_decap_8 FILLER_32_768 ();
 sg13g2_decap_8 FILLER_32_775 ();
 sg13g2_decap_8 FILLER_32_782 ();
 sg13g2_decap_8 FILLER_32_789 ();
 sg13g2_decap_8 FILLER_32_796 ();
 sg13g2_decap_8 FILLER_32_803 ();
 sg13g2_decap_8 FILLER_32_810 ();
 sg13g2_decap_8 FILLER_32_817 ();
 sg13g2_decap_8 FILLER_32_824 ();
 sg13g2_decap_8 FILLER_32_831 ();
 sg13g2_decap_8 FILLER_32_838 ();
 sg13g2_decap_8 FILLER_32_845 ();
 sg13g2_decap_8 FILLER_32_852 ();
 sg13g2_decap_8 FILLER_32_859 ();
 sg13g2_decap_8 FILLER_32_866 ();
 sg13g2_decap_8 FILLER_32_873 ();
 sg13g2_decap_8 FILLER_32_880 ();
 sg13g2_decap_8 FILLER_32_887 ();
 sg13g2_decap_8 FILLER_32_894 ();
 sg13g2_decap_8 FILLER_32_901 ();
 sg13g2_decap_8 FILLER_32_908 ();
 sg13g2_decap_8 FILLER_32_915 ();
 sg13g2_decap_8 FILLER_32_922 ();
 sg13g2_decap_8 FILLER_32_929 ();
 sg13g2_decap_8 FILLER_32_936 ();
 sg13g2_decap_8 FILLER_32_943 ();
 sg13g2_decap_8 FILLER_32_950 ();
 sg13g2_decap_8 FILLER_32_957 ();
 sg13g2_decap_8 FILLER_32_964 ();
 sg13g2_decap_8 FILLER_32_971 ();
 sg13g2_decap_8 FILLER_32_978 ();
 sg13g2_decap_8 FILLER_32_985 ();
 sg13g2_decap_8 FILLER_32_992 ();
 sg13g2_decap_8 FILLER_32_999 ();
 sg13g2_decap_8 FILLER_32_1006 ();
 sg13g2_decap_8 FILLER_32_1013 ();
 sg13g2_decap_8 FILLER_32_1020 ();
 sg13g2_fill_2 FILLER_32_1027 ();
 sg13g2_decap_8 FILLER_33_5 ();
 sg13g2_decap_8 FILLER_33_12 ();
 sg13g2_decap_8 FILLER_33_19 ();
 sg13g2_decap_8 FILLER_33_26 ();
 sg13g2_decap_8 FILLER_33_33 ();
 sg13g2_decap_8 FILLER_33_40 ();
 sg13g2_decap_8 FILLER_33_47 ();
 sg13g2_decap_8 FILLER_33_54 ();
 sg13g2_decap_8 FILLER_33_61 ();
 sg13g2_decap_8 FILLER_33_68 ();
 sg13g2_decap_8 FILLER_33_75 ();
 sg13g2_decap_8 FILLER_33_82 ();
 sg13g2_decap_8 FILLER_33_89 ();
 sg13g2_decap_8 FILLER_33_96 ();
 sg13g2_decap_8 FILLER_33_103 ();
 sg13g2_decap_8 FILLER_33_110 ();
 sg13g2_decap_8 FILLER_33_117 ();
 sg13g2_decap_8 FILLER_33_124 ();
 sg13g2_decap_8 FILLER_33_131 ();
 sg13g2_decap_8 FILLER_33_138 ();
 sg13g2_fill_2 FILLER_33_145 ();
 sg13g2_fill_1 FILLER_33_147 ();
 sg13g2_decap_8 FILLER_33_175 ();
 sg13g2_decap_8 FILLER_33_182 ();
 sg13g2_decap_8 FILLER_33_189 ();
 sg13g2_decap_8 FILLER_33_196 ();
 sg13g2_decap_8 FILLER_33_203 ();
 sg13g2_decap_8 FILLER_33_210 ();
 sg13g2_decap_8 FILLER_33_222 ();
 sg13g2_decap_8 FILLER_33_229 ();
 sg13g2_decap_8 FILLER_33_236 ();
 sg13g2_decap_8 FILLER_33_243 ();
 sg13g2_decap_8 FILLER_33_250 ();
 sg13g2_decap_4 FILLER_33_257 ();
 sg13g2_fill_1 FILLER_33_261 ();
 sg13g2_decap_4 FILLER_33_279 ();
 sg13g2_fill_2 FILLER_33_283 ();
 sg13g2_decap_8 FILLER_33_291 ();
 sg13g2_decap_8 FILLER_33_298 ();
 sg13g2_decap_8 FILLER_33_305 ();
 sg13g2_decap_8 FILLER_33_312 ();
 sg13g2_decap_8 FILLER_33_319 ();
 sg13g2_decap_8 FILLER_33_326 ();
 sg13g2_decap_8 FILLER_33_333 ();
 sg13g2_decap_8 FILLER_33_340 ();
 sg13g2_decap_4 FILLER_33_347 ();
 sg13g2_decap_8 FILLER_33_364 ();
 sg13g2_decap_8 FILLER_33_371 ();
 sg13g2_decap_8 FILLER_33_378 ();
 sg13g2_decap_8 FILLER_33_385 ();
 sg13g2_decap_8 FILLER_33_392 ();
 sg13g2_decap_4 FILLER_33_399 ();
 sg13g2_fill_2 FILLER_33_403 ();
 sg13g2_decap_8 FILLER_33_418 ();
 sg13g2_decap_8 FILLER_33_425 ();
 sg13g2_decap_8 FILLER_33_432 ();
 sg13g2_decap_8 FILLER_33_439 ();
 sg13g2_decap_8 FILLER_33_446 ();
 sg13g2_decap_8 FILLER_33_453 ();
 sg13g2_decap_8 FILLER_33_460 ();
 sg13g2_decap_8 FILLER_33_467 ();
 sg13g2_decap_8 FILLER_33_474 ();
 sg13g2_decap_8 FILLER_33_481 ();
 sg13g2_decap_8 FILLER_33_488 ();
 sg13g2_decap_8 FILLER_33_495 ();
 sg13g2_decap_8 FILLER_33_502 ();
 sg13g2_decap_8 FILLER_33_509 ();
 sg13g2_decap_8 FILLER_33_516 ();
 sg13g2_decap_8 FILLER_33_523 ();
 sg13g2_decap_8 FILLER_33_530 ();
 sg13g2_decap_8 FILLER_33_537 ();
 sg13g2_decap_8 FILLER_33_544 ();
 sg13g2_decap_8 FILLER_33_551 ();
 sg13g2_decap_8 FILLER_33_558 ();
 sg13g2_decap_8 FILLER_33_565 ();
 sg13g2_decap_8 FILLER_33_572 ();
 sg13g2_decap_8 FILLER_33_579 ();
 sg13g2_decap_8 FILLER_33_586 ();
 sg13g2_decap_8 FILLER_33_593 ();
 sg13g2_decap_8 FILLER_33_600 ();
 sg13g2_decap_8 FILLER_33_607 ();
 sg13g2_decap_8 FILLER_33_614 ();
 sg13g2_decap_8 FILLER_33_621 ();
 sg13g2_decap_8 FILLER_33_628 ();
 sg13g2_decap_8 FILLER_33_635 ();
 sg13g2_decap_8 FILLER_33_642 ();
 sg13g2_decap_8 FILLER_33_649 ();
 sg13g2_decap_8 FILLER_33_656 ();
 sg13g2_decap_8 FILLER_33_663 ();
 sg13g2_decap_8 FILLER_33_670 ();
 sg13g2_decap_8 FILLER_33_677 ();
 sg13g2_decap_8 FILLER_33_684 ();
 sg13g2_decap_8 FILLER_33_691 ();
 sg13g2_decap_8 FILLER_33_698 ();
 sg13g2_decap_8 FILLER_33_705 ();
 sg13g2_decap_8 FILLER_33_712 ();
 sg13g2_decap_8 FILLER_33_719 ();
 sg13g2_decap_8 FILLER_33_726 ();
 sg13g2_decap_8 FILLER_33_733 ();
 sg13g2_decap_8 FILLER_33_740 ();
 sg13g2_decap_8 FILLER_33_747 ();
 sg13g2_decap_8 FILLER_33_754 ();
 sg13g2_decap_8 FILLER_33_761 ();
 sg13g2_decap_8 FILLER_33_768 ();
 sg13g2_decap_8 FILLER_33_775 ();
 sg13g2_decap_8 FILLER_33_782 ();
 sg13g2_decap_8 FILLER_33_789 ();
 sg13g2_decap_8 FILLER_33_796 ();
 sg13g2_decap_8 FILLER_33_803 ();
 sg13g2_decap_8 FILLER_33_810 ();
 sg13g2_decap_8 FILLER_33_817 ();
 sg13g2_decap_8 FILLER_33_824 ();
 sg13g2_decap_8 FILLER_33_831 ();
 sg13g2_decap_8 FILLER_33_838 ();
 sg13g2_decap_8 FILLER_33_845 ();
 sg13g2_decap_8 FILLER_33_852 ();
 sg13g2_decap_8 FILLER_33_859 ();
 sg13g2_decap_8 FILLER_33_866 ();
 sg13g2_decap_8 FILLER_33_873 ();
 sg13g2_decap_8 FILLER_33_880 ();
 sg13g2_decap_8 FILLER_33_887 ();
 sg13g2_decap_8 FILLER_33_894 ();
 sg13g2_decap_8 FILLER_33_901 ();
 sg13g2_decap_8 FILLER_33_908 ();
 sg13g2_decap_8 FILLER_33_915 ();
 sg13g2_decap_8 FILLER_33_922 ();
 sg13g2_decap_8 FILLER_33_929 ();
 sg13g2_decap_8 FILLER_33_936 ();
 sg13g2_decap_8 FILLER_33_943 ();
 sg13g2_decap_8 FILLER_33_950 ();
 sg13g2_decap_8 FILLER_33_957 ();
 sg13g2_decap_8 FILLER_33_964 ();
 sg13g2_decap_8 FILLER_33_971 ();
 sg13g2_decap_8 FILLER_33_978 ();
 sg13g2_decap_8 FILLER_33_985 ();
 sg13g2_decap_8 FILLER_33_992 ();
 sg13g2_decap_8 FILLER_33_999 ();
 sg13g2_decap_8 FILLER_33_1006 ();
 sg13g2_decap_8 FILLER_33_1013 ();
 sg13g2_decap_8 FILLER_33_1020 ();
 sg13g2_fill_2 FILLER_33_1027 ();
 sg13g2_decap_8 FILLER_34_5 ();
 sg13g2_decap_8 FILLER_34_12 ();
 sg13g2_decap_8 FILLER_34_19 ();
 sg13g2_decap_8 FILLER_34_26 ();
 sg13g2_decap_8 FILLER_34_33 ();
 sg13g2_decap_8 FILLER_34_40 ();
 sg13g2_decap_8 FILLER_34_47 ();
 sg13g2_decap_8 FILLER_34_54 ();
 sg13g2_decap_8 FILLER_34_61 ();
 sg13g2_decap_8 FILLER_34_68 ();
 sg13g2_decap_8 FILLER_34_75 ();
 sg13g2_decap_8 FILLER_34_82 ();
 sg13g2_decap_8 FILLER_34_89 ();
 sg13g2_decap_8 FILLER_34_96 ();
 sg13g2_decap_8 FILLER_34_103 ();
 sg13g2_decap_8 FILLER_34_110 ();
 sg13g2_decap_8 FILLER_34_117 ();
 sg13g2_decap_8 FILLER_34_124 ();
 sg13g2_decap_8 FILLER_34_131 ();
 sg13g2_decap_8 FILLER_34_138 ();
 sg13g2_decap_8 FILLER_34_145 ();
 sg13g2_decap_8 FILLER_34_152 ();
 sg13g2_decap_8 FILLER_34_159 ();
 sg13g2_decap_8 FILLER_34_166 ();
 sg13g2_decap_8 FILLER_34_173 ();
 sg13g2_decap_8 FILLER_34_180 ();
 sg13g2_decap_8 FILLER_34_187 ();
 sg13g2_decap_4 FILLER_34_194 ();
 sg13g2_fill_2 FILLER_34_198 ();
 sg13g2_decap_8 FILLER_34_210 ();
 sg13g2_decap_8 FILLER_34_217 ();
 sg13g2_decap_8 FILLER_34_224 ();
 sg13g2_decap_8 FILLER_34_231 ();
 sg13g2_decap_8 FILLER_34_238 ();
 sg13g2_decap_8 FILLER_34_245 ();
 sg13g2_decap_8 FILLER_34_252 ();
 sg13g2_decap_8 FILLER_34_259 ();
 sg13g2_decap_8 FILLER_34_266 ();
 sg13g2_decap_8 FILLER_34_273 ();
 sg13g2_decap_8 FILLER_34_280 ();
 sg13g2_decap_8 FILLER_34_287 ();
 sg13g2_decap_4 FILLER_34_294 ();
 sg13g2_fill_2 FILLER_34_298 ();
 sg13g2_decap_8 FILLER_34_310 ();
 sg13g2_decap_8 FILLER_34_317 ();
 sg13g2_decap_8 FILLER_34_324 ();
 sg13g2_decap_8 FILLER_34_331 ();
 sg13g2_decap_8 FILLER_34_338 ();
 sg13g2_decap_8 FILLER_34_345 ();
 sg13g2_decap_4 FILLER_34_352 ();
 sg13g2_fill_1 FILLER_34_356 ();
 sg13g2_decap_8 FILLER_34_384 ();
 sg13g2_decap_8 FILLER_34_391 ();
 sg13g2_decap_8 FILLER_34_398 ();
 sg13g2_decap_8 FILLER_34_405 ();
 sg13g2_decap_8 FILLER_34_412 ();
 sg13g2_decap_8 FILLER_34_419 ();
 sg13g2_decap_8 FILLER_34_426 ();
 sg13g2_decap_8 FILLER_34_433 ();
 sg13g2_decap_8 FILLER_34_440 ();
 sg13g2_decap_8 FILLER_34_447 ();
 sg13g2_decap_8 FILLER_34_454 ();
 sg13g2_decap_8 FILLER_34_461 ();
 sg13g2_decap_8 FILLER_34_468 ();
 sg13g2_decap_8 FILLER_34_475 ();
 sg13g2_decap_8 FILLER_34_482 ();
 sg13g2_decap_8 FILLER_34_489 ();
 sg13g2_decap_8 FILLER_34_496 ();
 sg13g2_decap_8 FILLER_34_503 ();
 sg13g2_decap_8 FILLER_34_510 ();
 sg13g2_decap_8 FILLER_34_517 ();
 sg13g2_decap_8 FILLER_34_524 ();
 sg13g2_decap_8 FILLER_34_531 ();
 sg13g2_decap_8 FILLER_34_538 ();
 sg13g2_decap_8 FILLER_34_545 ();
 sg13g2_decap_8 FILLER_34_552 ();
 sg13g2_decap_8 FILLER_34_559 ();
 sg13g2_decap_8 FILLER_34_566 ();
 sg13g2_decap_8 FILLER_34_573 ();
 sg13g2_decap_8 FILLER_34_580 ();
 sg13g2_decap_8 FILLER_34_587 ();
 sg13g2_decap_8 FILLER_34_594 ();
 sg13g2_decap_8 FILLER_34_601 ();
 sg13g2_decap_8 FILLER_34_608 ();
 sg13g2_decap_8 FILLER_34_615 ();
 sg13g2_decap_8 FILLER_34_622 ();
 sg13g2_decap_8 FILLER_34_629 ();
 sg13g2_decap_8 FILLER_34_636 ();
 sg13g2_decap_8 FILLER_34_643 ();
 sg13g2_decap_8 FILLER_34_650 ();
 sg13g2_decap_8 FILLER_34_657 ();
 sg13g2_decap_8 FILLER_34_664 ();
 sg13g2_decap_8 FILLER_34_671 ();
 sg13g2_decap_8 FILLER_34_678 ();
 sg13g2_decap_8 FILLER_34_685 ();
 sg13g2_decap_8 FILLER_34_692 ();
 sg13g2_decap_8 FILLER_34_699 ();
 sg13g2_decap_8 FILLER_34_706 ();
 sg13g2_decap_8 FILLER_34_713 ();
 sg13g2_decap_8 FILLER_34_720 ();
 sg13g2_decap_8 FILLER_34_727 ();
 sg13g2_decap_8 FILLER_34_734 ();
 sg13g2_decap_8 FILLER_34_741 ();
 sg13g2_decap_8 FILLER_34_748 ();
 sg13g2_decap_8 FILLER_34_755 ();
 sg13g2_decap_8 FILLER_34_762 ();
 sg13g2_decap_8 FILLER_34_769 ();
 sg13g2_decap_8 FILLER_34_776 ();
 sg13g2_decap_8 FILLER_34_783 ();
 sg13g2_decap_8 FILLER_34_790 ();
 sg13g2_decap_8 FILLER_34_797 ();
 sg13g2_decap_8 FILLER_34_804 ();
 sg13g2_decap_8 FILLER_34_811 ();
 sg13g2_decap_8 FILLER_34_818 ();
 sg13g2_decap_8 FILLER_34_825 ();
 sg13g2_decap_8 FILLER_34_832 ();
 sg13g2_decap_8 FILLER_34_839 ();
 sg13g2_decap_8 FILLER_34_846 ();
 sg13g2_decap_8 FILLER_34_853 ();
 sg13g2_decap_8 FILLER_34_860 ();
 sg13g2_decap_8 FILLER_34_867 ();
 sg13g2_decap_8 FILLER_34_874 ();
 sg13g2_decap_8 FILLER_34_881 ();
 sg13g2_decap_8 FILLER_34_888 ();
 sg13g2_decap_8 FILLER_34_895 ();
 sg13g2_decap_8 FILLER_34_902 ();
 sg13g2_decap_8 FILLER_34_909 ();
 sg13g2_decap_8 FILLER_34_916 ();
 sg13g2_decap_8 FILLER_34_923 ();
 sg13g2_decap_8 FILLER_34_930 ();
 sg13g2_decap_8 FILLER_34_937 ();
 sg13g2_decap_8 FILLER_34_944 ();
 sg13g2_decap_8 FILLER_34_951 ();
 sg13g2_decap_8 FILLER_34_958 ();
 sg13g2_decap_8 FILLER_34_965 ();
 sg13g2_decap_8 FILLER_34_972 ();
 sg13g2_decap_8 FILLER_34_979 ();
 sg13g2_decap_8 FILLER_34_986 ();
 sg13g2_decap_8 FILLER_34_993 ();
 sg13g2_decap_8 FILLER_34_1000 ();
 sg13g2_decap_8 FILLER_34_1007 ();
 sg13g2_decap_8 FILLER_34_1014 ();
 sg13g2_decap_8 FILLER_34_1021 ();
 sg13g2_fill_1 FILLER_34_1028 ();
 sg13g2_decap_8 FILLER_35_5 ();
 sg13g2_decap_8 FILLER_35_12 ();
 sg13g2_decap_8 FILLER_35_19 ();
 sg13g2_decap_8 FILLER_35_26 ();
 sg13g2_decap_8 FILLER_35_33 ();
 sg13g2_decap_8 FILLER_35_40 ();
 sg13g2_decap_8 FILLER_35_47 ();
 sg13g2_decap_8 FILLER_35_54 ();
 sg13g2_decap_8 FILLER_35_61 ();
 sg13g2_decap_8 FILLER_35_68 ();
 sg13g2_decap_8 FILLER_35_75 ();
 sg13g2_decap_8 FILLER_35_82 ();
 sg13g2_decap_8 FILLER_35_89 ();
 sg13g2_decap_8 FILLER_35_96 ();
 sg13g2_decap_8 FILLER_35_103 ();
 sg13g2_decap_8 FILLER_35_110 ();
 sg13g2_decap_8 FILLER_35_117 ();
 sg13g2_decap_8 FILLER_35_124 ();
 sg13g2_decap_8 FILLER_35_131 ();
 sg13g2_decap_8 FILLER_35_138 ();
 sg13g2_decap_8 FILLER_35_145 ();
 sg13g2_decap_8 FILLER_35_152 ();
 sg13g2_decap_8 FILLER_35_159 ();
 sg13g2_decap_8 FILLER_35_166 ();
 sg13g2_decap_8 FILLER_35_173 ();
 sg13g2_fill_2 FILLER_35_180 ();
 sg13g2_decap_8 FILLER_35_192 ();
 sg13g2_fill_2 FILLER_35_199 ();
 sg13g2_fill_1 FILLER_35_201 ();
 sg13g2_decap_8 FILLER_35_207 ();
 sg13g2_decap_8 FILLER_35_214 ();
 sg13g2_decap_8 FILLER_35_221 ();
 sg13g2_decap_8 FILLER_35_228 ();
 sg13g2_fill_1 FILLER_35_235 ();
 sg13g2_decap_8 FILLER_35_241 ();
 sg13g2_decap_8 FILLER_35_248 ();
 sg13g2_decap_8 FILLER_35_255 ();
 sg13g2_decap_4 FILLER_35_262 ();
 sg13g2_fill_2 FILLER_35_266 ();
 sg13g2_decap_8 FILLER_35_278 ();
 sg13g2_decap_8 FILLER_35_285 ();
 sg13g2_decap_4 FILLER_35_292 ();
 sg13g2_fill_2 FILLER_35_296 ();
 sg13g2_decap_8 FILLER_35_304 ();
 sg13g2_decap_8 FILLER_35_311 ();
 sg13g2_decap_8 FILLER_35_318 ();
 sg13g2_decap_8 FILLER_35_325 ();
 sg13g2_decap_8 FILLER_35_332 ();
 sg13g2_decap_8 FILLER_35_339 ();
 sg13g2_decap_8 FILLER_35_346 ();
 sg13g2_decap_8 FILLER_35_353 ();
 sg13g2_decap_8 FILLER_35_360 ();
 sg13g2_decap_8 FILLER_35_367 ();
 sg13g2_decap_8 FILLER_35_374 ();
 sg13g2_decap_8 FILLER_35_381 ();
 sg13g2_decap_8 FILLER_35_388 ();
 sg13g2_decap_8 FILLER_35_395 ();
 sg13g2_decap_8 FILLER_35_402 ();
 sg13g2_decap_8 FILLER_35_409 ();
 sg13g2_decap_8 FILLER_35_416 ();
 sg13g2_decap_8 FILLER_35_423 ();
 sg13g2_decap_8 FILLER_35_430 ();
 sg13g2_decap_8 FILLER_35_437 ();
 sg13g2_decap_8 FILLER_35_444 ();
 sg13g2_decap_8 FILLER_35_451 ();
 sg13g2_decap_8 FILLER_35_458 ();
 sg13g2_decap_8 FILLER_35_465 ();
 sg13g2_decap_8 FILLER_35_472 ();
 sg13g2_decap_8 FILLER_35_479 ();
 sg13g2_decap_8 FILLER_35_486 ();
 sg13g2_decap_8 FILLER_35_493 ();
 sg13g2_decap_8 FILLER_35_500 ();
 sg13g2_decap_8 FILLER_35_507 ();
 sg13g2_decap_8 FILLER_35_514 ();
 sg13g2_decap_8 FILLER_35_521 ();
 sg13g2_decap_8 FILLER_35_528 ();
 sg13g2_decap_8 FILLER_35_535 ();
 sg13g2_decap_8 FILLER_35_542 ();
 sg13g2_decap_8 FILLER_35_549 ();
 sg13g2_decap_8 FILLER_35_556 ();
 sg13g2_decap_8 FILLER_35_563 ();
 sg13g2_decap_8 FILLER_35_570 ();
 sg13g2_decap_8 FILLER_35_577 ();
 sg13g2_decap_8 FILLER_35_584 ();
 sg13g2_decap_8 FILLER_35_591 ();
 sg13g2_decap_8 FILLER_35_598 ();
 sg13g2_decap_8 FILLER_35_605 ();
 sg13g2_decap_8 FILLER_35_612 ();
 sg13g2_decap_8 FILLER_35_619 ();
 sg13g2_decap_8 FILLER_35_626 ();
 sg13g2_decap_8 FILLER_35_633 ();
 sg13g2_decap_8 FILLER_35_640 ();
 sg13g2_decap_8 FILLER_35_647 ();
 sg13g2_decap_8 FILLER_35_654 ();
 sg13g2_decap_8 FILLER_35_661 ();
 sg13g2_decap_8 FILLER_35_668 ();
 sg13g2_decap_8 FILLER_35_675 ();
 sg13g2_decap_8 FILLER_35_682 ();
 sg13g2_decap_8 FILLER_35_689 ();
 sg13g2_decap_8 FILLER_35_696 ();
 sg13g2_decap_8 FILLER_35_703 ();
 sg13g2_decap_8 FILLER_35_710 ();
 sg13g2_decap_8 FILLER_35_717 ();
 sg13g2_decap_8 FILLER_35_724 ();
 sg13g2_decap_8 FILLER_35_731 ();
 sg13g2_decap_8 FILLER_35_738 ();
 sg13g2_decap_8 FILLER_35_745 ();
 sg13g2_decap_8 FILLER_35_752 ();
 sg13g2_decap_8 FILLER_35_759 ();
 sg13g2_decap_8 FILLER_35_766 ();
 sg13g2_decap_8 FILLER_35_773 ();
 sg13g2_decap_8 FILLER_35_780 ();
 sg13g2_decap_8 FILLER_35_787 ();
 sg13g2_decap_8 FILLER_35_794 ();
 sg13g2_decap_8 FILLER_35_801 ();
 sg13g2_decap_8 FILLER_35_808 ();
 sg13g2_decap_8 FILLER_35_815 ();
 sg13g2_decap_8 FILLER_35_822 ();
 sg13g2_decap_8 FILLER_35_829 ();
 sg13g2_decap_8 FILLER_35_836 ();
 sg13g2_decap_8 FILLER_35_843 ();
 sg13g2_decap_8 FILLER_35_850 ();
 sg13g2_decap_8 FILLER_35_857 ();
 sg13g2_decap_8 FILLER_35_864 ();
 sg13g2_decap_8 FILLER_35_871 ();
 sg13g2_decap_8 FILLER_35_878 ();
 sg13g2_decap_8 FILLER_35_885 ();
 sg13g2_decap_8 FILLER_35_892 ();
 sg13g2_decap_8 FILLER_35_899 ();
 sg13g2_decap_8 FILLER_35_906 ();
 sg13g2_decap_8 FILLER_35_913 ();
 sg13g2_decap_8 FILLER_35_920 ();
 sg13g2_decap_8 FILLER_35_927 ();
 sg13g2_decap_8 FILLER_35_934 ();
 sg13g2_decap_8 FILLER_35_941 ();
 sg13g2_decap_8 FILLER_35_948 ();
 sg13g2_decap_8 FILLER_35_955 ();
 sg13g2_decap_8 FILLER_35_962 ();
 sg13g2_decap_8 FILLER_35_969 ();
 sg13g2_decap_8 FILLER_35_976 ();
 sg13g2_decap_8 FILLER_35_983 ();
 sg13g2_decap_8 FILLER_35_990 ();
 sg13g2_decap_8 FILLER_35_997 ();
 sg13g2_decap_8 FILLER_35_1004 ();
 sg13g2_decap_8 FILLER_35_1011 ();
 sg13g2_decap_8 FILLER_35_1018 ();
 sg13g2_decap_4 FILLER_35_1025 ();
 sg13g2_decap_8 FILLER_36_5 ();
 sg13g2_decap_8 FILLER_36_12 ();
 sg13g2_decap_8 FILLER_36_19 ();
 sg13g2_decap_8 FILLER_36_26 ();
 sg13g2_decap_8 FILLER_36_33 ();
 sg13g2_decap_8 FILLER_36_40 ();
 sg13g2_decap_8 FILLER_36_47 ();
 sg13g2_decap_8 FILLER_36_54 ();
 sg13g2_decap_8 FILLER_36_61 ();
 sg13g2_decap_8 FILLER_36_68 ();
 sg13g2_decap_8 FILLER_36_75 ();
 sg13g2_decap_8 FILLER_36_82 ();
 sg13g2_decap_8 FILLER_36_89 ();
 sg13g2_decap_8 FILLER_36_96 ();
 sg13g2_decap_8 FILLER_36_103 ();
 sg13g2_decap_8 FILLER_36_110 ();
 sg13g2_decap_8 FILLER_36_117 ();
 sg13g2_decap_8 FILLER_36_124 ();
 sg13g2_decap_8 FILLER_36_131 ();
 sg13g2_decap_8 FILLER_36_138 ();
 sg13g2_decap_8 FILLER_36_145 ();
 sg13g2_decap_8 FILLER_36_152 ();
 sg13g2_decap_8 FILLER_36_159 ();
 sg13g2_decap_8 FILLER_36_166 ();
 sg13g2_decap_8 FILLER_36_173 ();
 sg13g2_decap_8 FILLER_36_180 ();
 sg13g2_decap_8 FILLER_36_187 ();
 sg13g2_decap_8 FILLER_36_194 ();
 sg13g2_decap_8 FILLER_36_201 ();
 sg13g2_decap_8 FILLER_36_208 ();
 sg13g2_decap_8 FILLER_36_215 ();
 sg13g2_fill_1 FILLER_36_222 ();
 sg13g2_decap_4 FILLER_36_230 ();
 sg13g2_fill_1 FILLER_36_234 ();
 sg13g2_decap_8 FILLER_36_240 ();
 sg13g2_decap_8 FILLER_36_247 ();
 sg13g2_decap_8 FILLER_36_254 ();
 sg13g2_decap_8 FILLER_36_261 ();
 sg13g2_decap_8 FILLER_36_268 ();
 sg13g2_decap_8 FILLER_36_275 ();
 sg13g2_decap_4 FILLER_36_282 ();
 sg13g2_fill_1 FILLER_36_292 ();
 sg13g2_decap_8 FILLER_36_305 ();
 sg13g2_decap_8 FILLER_36_312 ();
 sg13g2_decap_8 FILLER_36_319 ();
 sg13g2_decap_8 FILLER_36_326 ();
 sg13g2_decap_8 FILLER_36_333 ();
 sg13g2_decap_8 FILLER_36_340 ();
 sg13g2_decap_8 FILLER_36_347 ();
 sg13g2_decap_8 FILLER_36_354 ();
 sg13g2_decap_8 FILLER_36_361 ();
 sg13g2_decap_8 FILLER_36_368 ();
 sg13g2_decap_8 FILLER_36_375 ();
 sg13g2_decap_8 FILLER_36_382 ();
 sg13g2_decap_8 FILLER_36_389 ();
 sg13g2_decap_8 FILLER_36_396 ();
 sg13g2_decap_8 FILLER_36_403 ();
 sg13g2_decap_8 FILLER_36_410 ();
 sg13g2_decap_8 FILLER_36_417 ();
 sg13g2_decap_8 FILLER_36_424 ();
 sg13g2_decap_8 FILLER_36_431 ();
 sg13g2_decap_8 FILLER_36_438 ();
 sg13g2_decap_8 FILLER_36_445 ();
 sg13g2_decap_8 FILLER_36_452 ();
 sg13g2_decap_8 FILLER_36_459 ();
 sg13g2_decap_8 FILLER_36_466 ();
 sg13g2_decap_8 FILLER_36_473 ();
 sg13g2_decap_8 FILLER_36_480 ();
 sg13g2_decap_8 FILLER_36_487 ();
 sg13g2_decap_8 FILLER_36_494 ();
 sg13g2_decap_8 FILLER_36_501 ();
 sg13g2_decap_8 FILLER_36_508 ();
 sg13g2_decap_8 FILLER_36_515 ();
 sg13g2_decap_8 FILLER_36_522 ();
 sg13g2_decap_8 FILLER_36_529 ();
 sg13g2_decap_8 FILLER_36_536 ();
 sg13g2_decap_8 FILLER_36_543 ();
 sg13g2_decap_8 FILLER_36_550 ();
 sg13g2_decap_8 FILLER_36_557 ();
 sg13g2_decap_8 FILLER_36_564 ();
 sg13g2_decap_8 FILLER_36_571 ();
 sg13g2_decap_8 FILLER_36_578 ();
 sg13g2_decap_8 FILLER_36_585 ();
 sg13g2_decap_8 FILLER_36_592 ();
 sg13g2_decap_8 FILLER_36_599 ();
 sg13g2_decap_8 FILLER_36_606 ();
 sg13g2_decap_8 FILLER_36_613 ();
 sg13g2_decap_8 FILLER_36_620 ();
 sg13g2_decap_8 FILLER_36_627 ();
 sg13g2_decap_8 FILLER_36_634 ();
 sg13g2_decap_8 FILLER_36_641 ();
 sg13g2_decap_8 FILLER_36_648 ();
 sg13g2_decap_8 FILLER_36_655 ();
 sg13g2_decap_8 FILLER_36_662 ();
 sg13g2_decap_8 FILLER_36_669 ();
 sg13g2_decap_8 FILLER_36_676 ();
 sg13g2_decap_8 FILLER_36_683 ();
 sg13g2_decap_8 FILLER_36_690 ();
 sg13g2_decap_8 FILLER_36_697 ();
 sg13g2_decap_8 FILLER_36_704 ();
 sg13g2_decap_8 FILLER_36_711 ();
 sg13g2_decap_8 FILLER_36_718 ();
 sg13g2_decap_8 FILLER_36_725 ();
 sg13g2_decap_8 FILLER_36_732 ();
 sg13g2_decap_8 FILLER_36_739 ();
 sg13g2_decap_8 FILLER_36_746 ();
 sg13g2_decap_8 FILLER_36_753 ();
 sg13g2_decap_8 FILLER_36_760 ();
 sg13g2_decap_8 FILLER_36_767 ();
 sg13g2_decap_8 FILLER_36_774 ();
 sg13g2_decap_8 FILLER_36_781 ();
 sg13g2_decap_8 FILLER_36_788 ();
 sg13g2_decap_8 FILLER_36_795 ();
 sg13g2_decap_8 FILLER_36_802 ();
 sg13g2_decap_8 FILLER_36_809 ();
 sg13g2_decap_8 FILLER_36_816 ();
 sg13g2_decap_8 FILLER_36_823 ();
 sg13g2_decap_8 FILLER_36_830 ();
 sg13g2_decap_8 FILLER_36_837 ();
 sg13g2_decap_8 FILLER_36_844 ();
 sg13g2_decap_8 FILLER_36_851 ();
 sg13g2_decap_8 FILLER_36_858 ();
 sg13g2_decap_8 FILLER_36_865 ();
 sg13g2_decap_8 FILLER_36_872 ();
 sg13g2_decap_8 FILLER_36_879 ();
 sg13g2_decap_8 FILLER_36_886 ();
 sg13g2_decap_8 FILLER_36_893 ();
 sg13g2_decap_8 FILLER_36_900 ();
 sg13g2_decap_8 FILLER_36_907 ();
 sg13g2_decap_8 FILLER_36_914 ();
 sg13g2_decap_8 FILLER_36_921 ();
 sg13g2_decap_8 FILLER_36_928 ();
 sg13g2_decap_8 FILLER_36_935 ();
 sg13g2_decap_8 FILLER_36_942 ();
 sg13g2_decap_8 FILLER_36_949 ();
 sg13g2_decap_8 FILLER_36_956 ();
 sg13g2_decap_8 FILLER_36_963 ();
 sg13g2_decap_8 FILLER_36_970 ();
 sg13g2_decap_8 FILLER_36_977 ();
 sg13g2_decap_8 FILLER_36_984 ();
 sg13g2_decap_8 FILLER_36_991 ();
 sg13g2_decap_8 FILLER_36_998 ();
 sg13g2_decap_8 FILLER_36_1005 ();
 sg13g2_decap_8 FILLER_36_1012 ();
 sg13g2_decap_8 FILLER_36_1019 ();
 sg13g2_fill_2 FILLER_36_1026 ();
 sg13g2_fill_1 FILLER_36_1028 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_decap_4 FILLER_37_147 ();
 sg13g2_fill_2 FILLER_37_151 ();
 sg13g2_decap_8 FILLER_37_180 ();
 sg13g2_decap_8 FILLER_37_187 ();
 sg13g2_decap_8 FILLER_37_194 ();
 sg13g2_decap_8 FILLER_37_201 ();
 sg13g2_decap_8 FILLER_37_208 ();
 sg13g2_decap_8 FILLER_37_215 ();
 sg13g2_decap_8 FILLER_37_222 ();
 sg13g2_decap_8 FILLER_37_229 ();
 sg13g2_decap_8 FILLER_37_236 ();
 sg13g2_decap_8 FILLER_37_243 ();
 sg13g2_decap_8 FILLER_37_250 ();
 sg13g2_decap_8 FILLER_37_257 ();
 sg13g2_decap_8 FILLER_37_264 ();
 sg13g2_decap_8 FILLER_37_271 ();
 sg13g2_decap_8 FILLER_37_278 ();
 sg13g2_decap_8 FILLER_37_285 ();
 sg13g2_decap_8 FILLER_37_292 ();
 sg13g2_decap_8 FILLER_37_299 ();
 sg13g2_decap_8 FILLER_37_306 ();
 sg13g2_decap_4 FILLER_37_313 ();
 sg13g2_fill_1 FILLER_37_317 ();
 sg13g2_decap_8 FILLER_37_321 ();
 sg13g2_decap_8 FILLER_37_328 ();
 sg13g2_decap_8 FILLER_37_335 ();
 sg13g2_decap_8 FILLER_37_342 ();
 sg13g2_decap_8 FILLER_37_349 ();
 sg13g2_decap_8 FILLER_37_356 ();
 sg13g2_fill_1 FILLER_37_363 ();
 sg13g2_decap_8 FILLER_37_370 ();
 sg13g2_decap_8 FILLER_37_377 ();
 sg13g2_decap_8 FILLER_37_384 ();
 sg13g2_decap_8 FILLER_37_391 ();
 sg13g2_decap_8 FILLER_37_398 ();
 sg13g2_decap_8 FILLER_37_405 ();
 sg13g2_decap_8 FILLER_37_412 ();
 sg13g2_decap_8 FILLER_37_419 ();
 sg13g2_decap_8 FILLER_37_426 ();
 sg13g2_decap_8 FILLER_37_433 ();
 sg13g2_decap_8 FILLER_37_440 ();
 sg13g2_decap_8 FILLER_37_447 ();
 sg13g2_decap_8 FILLER_37_454 ();
 sg13g2_decap_8 FILLER_37_461 ();
 sg13g2_decap_8 FILLER_37_468 ();
 sg13g2_decap_8 FILLER_37_475 ();
 sg13g2_decap_8 FILLER_37_482 ();
 sg13g2_decap_8 FILLER_37_489 ();
 sg13g2_decap_8 FILLER_37_496 ();
 sg13g2_decap_8 FILLER_37_503 ();
 sg13g2_decap_8 FILLER_37_510 ();
 sg13g2_decap_8 FILLER_37_517 ();
 sg13g2_decap_8 FILLER_37_524 ();
 sg13g2_decap_8 FILLER_37_531 ();
 sg13g2_decap_8 FILLER_37_538 ();
 sg13g2_decap_8 FILLER_37_545 ();
 sg13g2_decap_8 FILLER_37_552 ();
 sg13g2_decap_8 FILLER_37_559 ();
 sg13g2_decap_8 FILLER_37_566 ();
 sg13g2_decap_8 FILLER_37_573 ();
 sg13g2_decap_8 FILLER_37_580 ();
 sg13g2_decap_8 FILLER_37_587 ();
 sg13g2_decap_8 FILLER_37_594 ();
 sg13g2_decap_8 FILLER_37_601 ();
 sg13g2_decap_8 FILLER_37_608 ();
 sg13g2_decap_8 FILLER_37_615 ();
 sg13g2_decap_8 FILLER_37_622 ();
 sg13g2_decap_8 FILLER_37_629 ();
 sg13g2_decap_8 FILLER_37_636 ();
 sg13g2_decap_8 FILLER_37_643 ();
 sg13g2_decap_8 FILLER_37_650 ();
 sg13g2_decap_8 FILLER_37_657 ();
 sg13g2_decap_8 FILLER_37_664 ();
 sg13g2_decap_8 FILLER_37_671 ();
 sg13g2_decap_8 FILLER_37_678 ();
 sg13g2_decap_8 FILLER_37_685 ();
 sg13g2_decap_8 FILLER_37_692 ();
 sg13g2_decap_8 FILLER_37_699 ();
 sg13g2_decap_8 FILLER_37_706 ();
 sg13g2_decap_8 FILLER_37_713 ();
 sg13g2_decap_8 FILLER_37_720 ();
 sg13g2_decap_8 FILLER_37_727 ();
 sg13g2_decap_8 FILLER_37_734 ();
 sg13g2_decap_8 FILLER_37_741 ();
 sg13g2_decap_8 FILLER_37_748 ();
 sg13g2_decap_8 FILLER_37_755 ();
 sg13g2_decap_8 FILLER_37_762 ();
 sg13g2_decap_8 FILLER_37_769 ();
 sg13g2_decap_8 FILLER_37_776 ();
 sg13g2_decap_8 FILLER_37_783 ();
 sg13g2_decap_8 FILLER_37_790 ();
 sg13g2_decap_8 FILLER_37_797 ();
 sg13g2_decap_8 FILLER_37_804 ();
 sg13g2_decap_8 FILLER_37_811 ();
 sg13g2_decap_8 FILLER_37_818 ();
 sg13g2_decap_8 FILLER_37_825 ();
 sg13g2_decap_8 FILLER_37_832 ();
 sg13g2_decap_8 FILLER_37_839 ();
 sg13g2_decap_8 FILLER_37_846 ();
 sg13g2_decap_8 FILLER_37_853 ();
 sg13g2_decap_8 FILLER_37_860 ();
 sg13g2_decap_8 FILLER_37_867 ();
 sg13g2_decap_8 FILLER_37_874 ();
 sg13g2_decap_8 FILLER_37_881 ();
 sg13g2_decap_8 FILLER_37_888 ();
 sg13g2_decap_8 FILLER_37_895 ();
 sg13g2_decap_8 FILLER_37_902 ();
 sg13g2_decap_8 FILLER_37_909 ();
 sg13g2_decap_8 FILLER_37_916 ();
 sg13g2_decap_8 FILLER_37_923 ();
 sg13g2_decap_8 FILLER_37_930 ();
 sg13g2_decap_8 FILLER_37_937 ();
 sg13g2_decap_8 FILLER_37_944 ();
 sg13g2_decap_8 FILLER_37_951 ();
 sg13g2_decap_8 FILLER_37_958 ();
 sg13g2_decap_8 FILLER_37_965 ();
 sg13g2_decap_8 FILLER_37_972 ();
 sg13g2_decap_8 FILLER_37_979 ();
 sg13g2_decap_8 FILLER_37_986 ();
 sg13g2_decap_8 FILLER_37_993 ();
 sg13g2_decap_8 FILLER_37_1000 ();
 sg13g2_decap_8 FILLER_37_1007 ();
 sg13g2_decap_8 FILLER_37_1014 ();
 sg13g2_decap_8 FILLER_37_1021 ();
 sg13g2_fill_1 FILLER_37_1028 ();
 sg13g2_decap_8 FILLER_38_4 ();
 sg13g2_decap_8 FILLER_38_11 ();
 sg13g2_decap_8 FILLER_38_18 ();
 sg13g2_decap_8 FILLER_38_25 ();
 sg13g2_decap_8 FILLER_38_32 ();
 sg13g2_decap_8 FILLER_38_39 ();
 sg13g2_decap_8 FILLER_38_46 ();
 sg13g2_decap_8 FILLER_38_53 ();
 sg13g2_decap_8 FILLER_38_60 ();
 sg13g2_decap_8 FILLER_38_67 ();
 sg13g2_decap_8 FILLER_38_74 ();
 sg13g2_decap_8 FILLER_38_81 ();
 sg13g2_decap_8 FILLER_38_88 ();
 sg13g2_decap_8 FILLER_38_95 ();
 sg13g2_decap_8 FILLER_38_102 ();
 sg13g2_decap_8 FILLER_38_109 ();
 sg13g2_decap_8 FILLER_38_116 ();
 sg13g2_decap_8 FILLER_38_123 ();
 sg13g2_decap_8 FILLER_38_130 ();
 sg13g2_decap_8 FILLER_38_137 ();
 sg13g2_decap_8 FILLER_38_144 ();
 sg13g2_decap_8 FILLER_38_151 ();
 sg13g2_decap_8 FILLER_38_158 ();
 sg13g2_decap_8 FILLER_38_165 ();
 sg13g2_decap_8 FILLER_38_172 ();
 sg13g2_decap_8 FILLER_38_179 ();
 sg13g2_decap_8 FILLER_38_186 ();
 sg13g2_decap_8 FILLER_38_193 ();
 sg13g2_decap_8 FILLER_38_200 ();
 sg13g2_decap_8 FILLER_38_207 ();
 sg13g2_decap_8 FILLER_38_214 ();
 sg13g2_decap_8 FILLER_38_221 ();
 sg13g2_decap_8 FILLER_38_228 ();
 sg13g2_decap_8 FILLER_38_235 ();
 sg13g2_decap_8 FILLER_38_242 ();
 sg13g2_decap_8 FILLER_38_249 ();
 sg13g2_decap_8 FILLER_38_256 ();
 sg13g2_decap_8 FILLER_38_263 ();
 sg13g2_decap_8 FILLER_38_270 ();
 sg13g2_decap_8 FILLER_38_277 ();
 sg13g2_decap_8 FILLER_38_284 ();
 sg13g2_decap_8 FILLER_38_291 ();
 sg13g2_decap_8 FILLER_38_298 ();
 sg13g2_decap_8 FILLER_38_305 ();
 sg13g2_decap_8 FILLER_38_312 ();
 sg13g2_decap_8 FILLER_38_319 ();
 sg13g2_decap_8 FILLER_38_326 ();
 sg13g2_decap_8 FILLER_38_333 ();
 sg13g2_decap_8 FILLER_38_340 ();
 sg13g2_decap_8 FILLER_38_347 ();
 sg13g2_decap_8 FILLER_38_354 ();
 sg13g2_decap_8 FILLER_38_361 ();
 sg13g2_decap_4 FILLER_38_368 ();
 sg13g2_fill_1 FILLER_38_372 ();
 sg13g2_decap_8 FILLER_38_379 ();
 sg13g2_decap_8 FILLER_38_386 ();
 sg13g2_decap_8 FILLER_38_393 ();
 sg13g2_decap_8 FILLER_38_400 ();
 sg13g2_decap_8 FILLER_38_407 ();
 sg13g2_decap_8 FILLER_38_414 ();
 sg13g2_decap_8 FILLER_38_421 ();
 sg13g2_decap_8 FILLER_38_428 ();
 sg13g2_decap_8 FILLER_38_435 ();
 sg13g2_decap_8 FILLER_38_442 ();
 sg13g2_decap_8 FILLER_38_449 ();
 sg13g2_decap_8 FILLER_38_456 ();
 sg13g2_decap_8 FILLER_38_463 ();
 sg13g2_decap_8 FILLER_38_470 ();
 sg13g2_decap_8 FILLER_38_477 ();
 sg13g2_decap_8 FILLER_38_484 ();
 sg13g2_decap_8 FILLER_38_491 ();
 sg13g2_decap_8 FILLER_38_498 ();
 sg13g2_decap_8 FILLER_38_505 ();
 sg13g2_decap_8 FILLER_38_512 ();
 sg13g2_decap_8 FILLER_38_519 ();
 sg13g2_decap_8 FILLER_38_526 ();
 sg13g2_decap_8 FILLER_38_533 ();
 sg13g2_decap_8 FILLER_38_540 ();
 sg13g2_decap_8 FILLER_38_547 ();
 sg13g2_decap_8 FILLER_38_554 ();
 sg13g2_decap_8 FILLER_38_561 ();
 sg13g2_decap_8 FILLER_38_568 ();
 sg13g2_decap_8 FILLER_38_575 ();
 sg13g2_decap_8 FILLER_38_582 ();
 sg13g2_decap_8 FILLER_38_589 ();
 sg13g2_decap_8 FILLER_38_596 ();
 sg13g2_decap_8 FILLER_38_603 ();
 sg13g2_decap_8 FILLER_38_610 ();
 sg13g2_decap_8 FILLER_38_617 ();
 sg13g2_decap_8 FILLER_38_624 ();
 sg13g2_decap_8 FILLER_38_631 ();
 sg13g2_decap_8 FILLER_38_638 ();
 sg13g2_decap_8 FILLER_38_645 ();
 sg13g2_decap_8 FILLER_38_652 ();
 sg13g2_decap_8 FILLER_38_659 ();
 sg13g2_decap_8 FILLER_38_666 ();
 sg13g2_decap_8 FILLER_38_673 ();
 sg13g2_decap_8 FILLER_38_680 ();
 sg13g2_decap_8 FILLER_38_687 ();
 sg13g2_decap_8 FILLER_38_694 ();
 sg13g2_decap_8 FILLER_38_701 ();
 sg13g2_decap_8 FILLER_38_708 ();
 sg13g2_decap_8 FILLER_38_715 ();
 sg13g2_decap_8 FILLER_38_722 ();
 sg13g2_decap_8 FILLER_38_729 ();
 sg13g2_decap_8 FILLER_38_736 ();
 sg13g2_decap_8 FILLER_38_743 ();
 sg13g2_decap_8 FILLER_38_750 ();
 sg13g2_decap_8 FILLER_38_757 ();
 sg13g2_decap_8 FILLER_38_764 ();
 sg13g2_decap_8 FILLER_38_771 ();
 sg13g2_decap_8 FILLER_38_778 ();
 sg13g2_decap_8 FILLER_38_785 ();
 sg13g2_decap_8 FILLER_38_792 ();
 sg13g2_decap_8 FILLER_38_799 ();
 sg13g2_decap_8 FILLER_38_806 ();
 sg13g2_decap_8 FILLER_38_813 ();
 sg13g2_decap_8 FILLER_38_820 ();
 sg13g2_decap_8 FILLER_38_827 ();
 sg13g2_decap_8 FILLER_38_834 ();
 sg13g2_decap_8 FILLER_38_841 ();
 sg13g2_decap_8 FILLER_38_848 ();
 sg13g2_decap_8 FILLER_38_855 ();
 sg13g2_decap_8 FILLER_38_862 ();
 sg13g2_decap_8 FILLER_38_869 ();
 sg13g2_decap_8 FILLER_38_876 ();
 sg13g2_decap_8 FILLER_38_883 ();
 sg13g2_decap_8 FILLER_38_890 ();
 sg13g2_decap_8 FILLER_38_897 ();
 sg13g2_decap_8 FILLER_38_904 ();
 sg13g2_decap_8 FILLER_38_911 ();
 sg13g2_decap_8 FILLER_38_918 ();
 sg13g2_decap_8 FILLER_38_925 ();
 sg13g2_decap_8 FILLER_38_932 ();
 sg13g2_decap_8 FILLER_38_939 ();
 sg13g2_decap_8 FILLER_38_946 ();
 sg13g2_decap_8 FILLER_38_953 ();
 sg13g2_decap_8 FILLER_38_960 ();
 sg13g2_decap_8 FILLER_38_967 ();
 sg13g2_decap_8 FILLER_38_974 ();
 sg13g2_decap_8 FILLER_38_981 ();
 sg13g2_decap_8 FILLER_38_988 ();
 sg13g2_decap_8 FILLER_38_995 ();
 sg13g2_decap_8 FILLER_38_1002 ();
 sg13g2_decap_8 FILLER_38_1009 ();
 sg13g2_decap_8 FILLER_38_1016 ();
 sg13g2_decap_4 FILLER_38_1023 ();
 sg13g2_fill_2 FILLER_38_1027 ();
 sg13g2_decap_8 FILLER_39_4 ();
 sg13g2_decap_8 FILLER_39_11 ();
 sg13g2_decap_8 FILLER_39_18 ();
 sg13g2_decap_8 FILLER_39_25 ();
 sg13g2_decap_8 FILLER_39_32 ();
 sg13g2_decap_8 FILLER_39_39 ();
 sg13g2_decap_8 FILLER_39_46 ();
 sg13g2_decap_8 FILLER_39_53 ();
 sg13g2_decap_8 FILLER_39_60 ();
 sg13g2_decap_8 FILLER_39_67 ();
 sg13g2_decap_8 FILLER_39_74 ();
 sg13g2_decap_8 FILLER_39_81 ();
 sg13g2_decap_8 FILLER_39_88 ();
 sg13g2_decap_8 FILLER_39_95 ();
 sg13g2_decap_8 FILLER_39_102 ();
 sg13g2_decap_8 FILLER_39_109 ();
 sg13g2_decap_8 FILLER_39_116 ();
 sg13g2_decap_8 FILLER_39_123 ();
 sg13g2_decap_8 FILLER_39_130 ();
 sg13g2_decap_8 FILLER_39_137 ();
 sg13g2_decap_8 FILLER_39_144 ();
 sg13g2_decap_8 FILLER_39_151 ();
 sg13g2_decap_8 FILLER_39_158 ();
 sg13g2_decap_8 FILLER_39_165 ();
 sg13g2_decap_8 FILLER_39_172 ();
 sg13g2_decap_8 FILLER_39_179 ();
 sg13g2_decap_8 FILLER_39_186 ();
 sg13g2_decap_8 FILLER_39_193 ();
 sg13g2_decap_8 FILLER_39_200 ();
 sg13g2_decap_8 FILLER_39_207 ();
 sg13g2_decap_8 FILLER_39_214 ();
 sg13g2_decap_8 FILLER_39_221 ();
 sg13g2_decap_8 FILLER_39_228 ();
 sg13g2_decap_8 FILLER_39_235 ();
 sg13g2_decap_8 FILLER_39_242 ();
 sg13g2_decap_8 FILLER_39_249 ();
 sg13g2_decap_8 FILLER_39_256 ();
 sg13g2_decap_8 FILLER_39_263 ();
 sg13g2_decap_8 FILLER_39_270 ();
 sg13g2_decap_8 FILLER_39_283 ();
 sg13g2_decap_8 FILLER_39_290 ();
 sg13g2_decap_8 FILLER_39_297 ();
 sg13g2_decap_8 FILLER_39_304 ();
 sg13g2_decap_8 FILLER_39_311 ();
 sg13g2_decap_8 FILLER_39_318 ();
 sg13g2_decap_8 FILLER_39_325 ();
 sg13g2_fill_2 FILLER_39_332 ();
 sg13g2_decap_8 FILLER_39_361 ();
 sg13g2_decap_8 FILLER_39_368 ();
 sg13g2_decap_8 FILLER_39_375 ();
 sg13g2_decap_8 FILLER_39_382 ();
 sg13g2_decap_8 FILLER_39_389 ();
 sg13g2_decap_8 FILLER_39_396 ();
 sg13g2_decap_8 FILLER_39_403 ();
 sg13g2_decap_8 FILLER_39_410 ();
 sg13g2_decap_8 FILLER_39_417 ();
 sg13g2_decap_8 FILLER_39_424 ();
 sg13g2_decap_8 FILLER_39_431 ();
 sg13g2_decap_8 FILLER_39_438 ();
 sg13g2_decap_8 FILLER_39_445 ();
 sg13g2_decap_8 FILLER_39_452 ();
 sg13g2_decap_8 FILLER_39_459 ();
 sg13g2_decap_8 FILLER_39_466 ();
 sg13g2_decap_8 FILLER_39_473 ();
 sg13g2_decap_8 FILLER_39_480 ();
 sg13g2_decap_8 FILLER_39_487 ();
 sg13g2_decap_8 FILLER_39_494 ();
 sg13g2_decap_8 FILLER_39_501 ();
 sg13g2_decap_8 FILLER_39_508 ();
 sg13g2_decap_8 FILLER_39_515 ();
 sg13g2_decap_8 FILLER_39_522 ();
 sg13g2_decap_8 FILLER_39_529 ();
 sg13g2_decap_8 FILLER_39_536 ();
 sg13g2_decap_8 FILLER_39_543 ();
 sg13g2_decap_8 FILLER_39_550 ();
 sg13g2_decap_8 FILLER_39_557 ();
 sg13g2_decap_8 FILLER_39_564 ();
 sg13g2_decap_8 FILLER_39_571 ();
 sg13g2_decap_8 FILLER_39_578 ();
 sg13g2_decap_8 FILLER_39_585 ();
 sg13g2_decap_8 FILLER_39_592 ();
 sg13g2_decap_8 FILLER_39_599 ();
 sg13g2_decap_8 FILLER_39_606 ();
 sg13g2_decap_8 FILLER_39_613 ();
 sg13g2_decap_8 FILLER_39_620 ();
 sg13g2_decap_8 FILLER_39_627 ();
 sg13g2_decap_8 FILLER_39_634 ();
 sg13g2_decap_8 FILLER_39_641 ();
 sg13g2_decap_8 FILLER_39_648 ();
 sg13g2_decap_8 FILLER_39_655 ();
 sg13g2_decap_8 FILLER_39_662 ();
 sg13g2_decap_8 FILLER_39_669 ();
 sg13g2_decap_8 FILLER_39_676 ();
 sg13g2_decap_8 FILLER_39_683 ();
 sg13g2_decap_8 FILLER_39_690 ();
 sg13g2_decap_8 FILLER_39_697 ();
 sg13g2_decap_8 FILLER_39_704 ();
 sg13g2_decap_8 FILLER_39_711 ();
 sg13g2_decap_8 FILLER_39_718 ();
 sg13g2_decap_8 FILLER_39_725 ();
 sg13g2_decap_8 FILLER_39_732 ();
 sg13g2_decap_8 FILLER_39_739 ();
 sg13g2_decap_8 FILLER_39_746 ();
 sg13g2_decap_8 FILLER_39_753 ();
 sg13g2_decap_8 FILLER_39_760 ();
 sg13g2_decap_8 FILLER_39_767 ();
 sg13g2_decap_8 FILLER_39_774 ();
 sg13g2_decap_8 FILLER_39_781 ();
 sg13g2_decap_8 FILLER_39_788 ();
 sg13g2_decap_8 FILLER_39_795 ();
 sg13g2_decap_8 FILLER_39_802 ();
 sg13g2_decap_8 FILLER_39_809 ();
 sg13g2_decap_8 FILLER_39_816 ();
 sg13g2_decap_8 FILLER_39_823 ();
 sg13g2_decap_8 FILLER_39_830 ();
 sg13g2_decap_8 FILLER_39_837 ();
 sg13g2_decap_8 FILLER_39_844 ();
 sg13g2_decap_8 FILLER_39_851 ();
 sg13g2_decap_8 FILLER_39_858 ();
 sg13g2_decap_8 FILLER_39_865 ();
 sg13g2_decap_8 FILLER_39_872 ();
 sg13g2_decap_8 FILLER_39_879 ();
 sg13g2_decap_8 FILLER_39_886 ();
 sg13g2_decap_8 FILLER_39_893 ();
 sg13g2_decap_8 FILLER_39_900 ();
 sg13g2_decap_8 FILLER_39_907 ();
 sg13g2_decap_8 FILLER_39_914 ();
 sg13g2_decap_8 FILLER_39_921 ();
 sg13g2_decap_8 FILLER_39_928 ();
 sg13g2_decap_8 FILLER_39_935 ();
 sg13g2_decap_8 FILLER_39_942 ();
 sg13g2_decap_8 FILLER_39_949 ();
 sg13g2_decap_8 FILLER_39_956 ();
 sg13g2_decap_8 FILLER_39_963 ();
 sg13g2_decap_8 FILLER_39_970 ();
 sg13g2_decap_8 FILLER_39_977 ();
 sg13g2_decap_8 FILLER_39_984 ();
 sg13g2_decap_8 FILLER_39_991 ();
 sg13g2_decap_8 FILLER_39_998 ();
 sg13g2_decap_8 FILLER_39_1005 ();
 sg13g2_decap_8 FILLER_39_1012 ();
 sg13g2_decap_8 FILLER_39_1019 ();
 sg13g2_fill_2 FILLER_39_1026 ();
 sg13g2_fill_1 FILLER_39_1028 ();
 sg13g2_decap_8 FILLER_40_4 ();
 sg13g2_decap_8 FILLER_40_11 ();
 sg13g2_decap_8 FILLER_40_18 ();
 sg13g2_decap_8 FILLER_40_25 ();
 sg13g2_decap_8 FILLER_40_32 ();
 sg13g2_decap_8 FILLER_40_39 ();
 sg13g2_decap_8 FILLER_40_46 ();
 sg13g2_decap_8 FILLER_40_53 ();
 sg13g2_decap_8 FILLER_40_60 ();
 sg13g2_decap_8 FILLER_40_67 ();
 sg13g2_decap_8 FILLER_40_74 ();
 sg13g2_decap_8 FILLER_40_81 ();
 sg13g2_decap_8 FILLER_40_88 ();
 sg13g2_decap_8 FILLER_40_95 ();
 sg13g2_decap_8 FILLER_40_102 ();
 sg13g2_decap_8 FILLER_40_109 ();
 sg13g2_decap_8 FILLER_40_116 ();
 sg13g2_decap_8 FILLER_40_123 ();
 sg13g2_decap_8 FILLER_40_130 ();
 sg13g2_decap_8 FILLER_40_137 ();
 sg13g2_decap_8 FILLER_40_144 ();
 sg13g2_decap_8 FILLER_40_151 ();
 sg13g2_decap_8 FILLER_40_158 ();
 sg13g2_decap_8 FILLER_40_165 ();
 sg13g2_decap_8 FILLER_40_172 ();
 sg13g2_decap_8 FILLER_40_179 ();
 sg13g2_decap_8 FILLER_40_186 ();
 sg13g2_decap_8 FILLER_40_193 ();
 sg13g2_decap_8 FILLER_40_200 ();
 sg13g2_decap_8 FILLER_40_207 ();
 sg13g2_fill_2 FILLER_40_214 ();
 sg13g2_decap_8 FILLER_40_243 ();
 sg13g2_decap_8 FILLER_40_250 ();
 sg13g2_decap_8 FILLER_40_257 ();
 sg13g2_decap_8 FILLER_40_264 ();
 sg13g2_fill_1 FILLER_40_271 ();
 sg13g2_decap_8 FILLER_40_299 ();
 sg13g2_decap_8 FILLER_40_306 ();
 sg13g2_decap_8 FILLER_40_313 ();
 sg13g2_decap_8 FILLER_40_320 ();
 sg13g2_decap_8 FILLER_40_327 ();
 sg13g2_decap_8 FILLER_40_334 ();
 sg13g2_decap_8 FILLER_40_341 ();
 sg13g2_decap_8 FILLER_40_348 ();
 sg13g2_decap_8 FILLER_40_355 ();
 sg13g2_decap_8 FILLER_40_362 ();
 sg13g2_decap_8 FILLER_40_369 ();
 sg13g2_decap_8 FILLER_40_376 ();
 sg13g2_decap_8 FILLER_40_383 ();
 sg13g2_decap_8 FILLER_40_390 ();
 sg13g2_decap_8 FILLER_40_397 ();
 sg13g2_decap_8 FILLER_40_404 ();
 sg13g2_decap_8 FILLER_40_411 ();
 sg13g2_decap_8 FILLER_40_418 ();
 sg13g2_decap_8 FILLER_40_425 ();
 sg13g2_decap_8 FILLER_40_432 ();
 sg13g2_decap_8 FILLER_40_439 ();
 sg13g2_decap_8 FILLER_40_446 ();
 sg13g2_decap_8 FILLER_40_453 ();
 sg13g2_decap_8 FILLER_40_460 ();
 sg13g2_decap_8 FILLER_40_467 ();
 sg13g2_decap_8 FILLER_40_474 ();
 sg13g2_decap_8 FILLER_40_481 ();
 sg13g2_decap_8 FILLER_40_488 ();
 sg13g2_decap_8 FILLER_40_495 ();
 sg13g2_decap_8 FILLER_40_502 ();
 sg13g2_decap_8 FILLER_40_509 ();
 sg13g2_decap_8 FILLER_40_516 ();
 sg13g2_decap_8 FILLER_40_523 ();
 sg13g2_decap_8 FILLER_40_530 ();
 sg13g2_decap_8 FILLER_40_537 ();
 sg13g2_decap_8 FILLER_40_544 ();
 sg13g2_decap_8 FILLER_40_551 ();
 sg13g2_decap_8 FILLER_40_558 ();
 sg13g2_decap_8 FILLER_40_565 ();
 sg13g2_decap_8 FILLER_40_572 ();
 sg13g2_decap_8 FILLER_40_579 ();
 sg13g2_decap_8 FILLER_40_586 ();
 sg13g2_decap_8 FILLER_40_593 ();
 sg13g2_decap_8 FILLER_40_600 ();
 sg13g2_decap_8 FILLER_40_607 ();
 sg13g2_decap_8 FILLER_40_614 ();
 sg13g2_decap_8 FILLER_40_621 ();
 sg13g2_decap_8 FILLER_40_628 ();
 sg13g2_decap_8 FILLER_40_635 ();
 sg13g2_decap_8 FILLER_40_642 ();
 sg13g2_decap_8 FILLER_40_649 ();
 sg13g2_decap_8 FILLER_40_656 ();
 sg13g2_decap_8 FILLER_40_663 ();
 sg13g2_decap_8 FILLER_40_670 ();
 sg13g2_decap_8 FILLER_40_677 ();
 sg13g2_decap_8 FILLER_40_684 ();
 sg13g2_decap_8 FILLER_40_691 ();
 sg13g2_decap_8 FILLER_40_698 ();
 sg13g2_decap_8 FILLER_40_705 ();
 sg13g2_decap_8 FILLER_40_712 ();
 sg13g2_decap_8 FILLER_40_719 ();
 sg13g2_decap_8 FILLER_40_726 ();
 sg13g2_decap_8 FILLER_40_733 ();
 sg13g2_decap_8 FILLER_40_740 ();
 sg13g2_decap_8 FILLER_40_747 ();
 sg13g2_decap_8 FILLER_40_754 ();
 sg13g2_decap_8 FILLER_40_761 ();
 sg13g2_decap_8 FILLER_40_768 ();
 sg13g2_decap_8 FILLER_40_775 ();
 sg13g2_decap_8 FILLER_40_782 ();
 sg13g2_decap_8 FILLER_40_789 ();
 sg13g2_decap_8 FILLER_40_796 ();
 sg13g2_decap_8 FILLER_40_803 ();
 sg13g2_decap_8 FILLER_40_810 ();
 sg13g2_decap_8 FILLER_40_817 ();
 sg13g2_decap_8 FILLER_40_824 ();
 sg13g2_decap_8 FILLER_40_831 ();
 sg13g2_decap_8 FILLER_40_838 ();
 sg13g2_decap_8 FILLER_40_845 ();
 sg13g2_decap_8 FILLER_40_852 ();
 sg13g2_decap_8 FILLER_40_859 ();
 sg13g2_decap_8 FILLER_40_866 ();
 sg13g2_decap_8 FILLER_40_873 ();
 sg13g2_decap_8 FILLER_40_880 ();
 sg13g2_decap_8 FILLER_40_887 ();
 sg13g2_decap_8 FILLER_40_894 ();
 sg13g2_decap_8 FILLER_40_901 ();
 sg13g2_decap_8 FILLER_40_908 ();
 sg13g2_decap_8 FILLER_40_915 ();
 sg13g2_decap_8 FILLER_40_922 ();
 sg13g2_decap_8 FILLER_40_929 ();
 sg13g2_decap_8 FILLER_40_936 ();
 sg13g2_decap_8 FILLER_40_943 ();
 sg13g2_decap_8 FILLER_40_950 ();
 sg13g2_decap_8 FILLER_40_957 ();
 sg13g2_decap_8 FILLER_40_964 ();
 sg13g2_decap_8 FILLER_40_971 ();
 sg13g2_decap_8 FILLER_40_978 ();
 sg13g2_decap_8 FILLER_40_985 ();
 sg13g2_decap_8 FILLER_40_992 ();
 sg13g2_decap_8 FILLER_40_999 ();
 sg13g2_decap_8 FILLER_40_1006 ();
 sg13g2_decap_8 FILLER_40_1013 ();
 sg13g2_decap_8 FILLER_40_1020 ();
 sg13g2_fill_2 FILLER_40_1027 ();
 sg13g2_decap_8 FILLER_41_4 ();
 sg13g2_decap_8 FILLER_41_11 ();
 sg13g2_decap_8 FILLER_41_18 ();
 sg13g2_decap_8 FILLER_41_25 ();
 sg13g2_decap_8 FILLER_41_32 ();
 sg13g2_decap_8 FILLER_41_39 ();
 sg13g2_decap_8 FILLER_41_46 ();
 sg13g2_decap_8 FILLER_41_53 ();
 sg13g2_decap_8 FILLER_41_60 ();
 sg13g2_decap_8 FILLER_41_67 ();
 sg13g2_decap_8 FILLER_41_74 ();
 sg13g2_decap_8 FILLER_41_81 ();
 sg13g2_decap_8 FILLER_41_88 ();
 sg13g2_decap_8 FILLER_41_95 ();
 sg13g2_decap_8 FILLER_41_102 ();
 sg13g2_decap_8 FILLER_41_109 ();
 sg13g2_decap_8 FILLER_41_116 ();
 sg13g2_decap_8 FILLER_41_123 ();
 sg13g2_decap_8 FILLER_41_130 ();
 sg13g2_decap_8 FILLER_41_137 ();
 sg13g2_decap_8 FILLER_41_144 ();
 sg13g2_decap_8 FILLER_41_151 ();
 sg13g2_decap_8 FILLER_41_158 ();
 sg13g2_decap_8 FILLER_41_165 ();
 sg13g2_decap_8 FILLER_41_172 ();
 sg13g2_decap_8 FILLER_41_179 ();
 sg13g2_decap_8 FILLER_41_186 ();
 sg13g2_decap_8 FILLER_41_193 ();
 sg13g2_decap_8 FILLER_41_200 ();
 sg13g2_decap_8 FILLER_41_207 ();
 sg13g2_decap_8 FILLER_41_214 ();
 sg13g2_decap_8 FILLER_41_221 ();
 sg13g2_decap_8 FILLER_41_228 ();
 sg13g2_decap_8 FILLER_41_235 ();
 sg13g2_decap_8 FILLER_41_242 ();
 sg13g2_decap_8 FILLER_41_249 ();
 sg13g2_decap_8 FILLER_41_256 ();
 sg13g2_decap_8 FILLER_41_263 ();
 sg13g2_decap_8 FILLER_41_270 ();
 sg13g2_fill_2 FILLER_41_277 ();
 sg13g2_decap_8 FILLER_41_285 ();
 sg13g2_decap_8 FILLER_41_292 ();
 sg13g2_decap_8 FILLER_41_299 ();
 sg13g2_decap_8 FILLER_41_306 ();
 sg13g2_decap_8 FILLER_41_313 ();
 sg13g2_decap_8 FILLER_41_320 ();
 sg13g2_decap_8 FILLER_41_327 ();
 sg13g2_decap_8 FILLER_41_334 ();
 sg13g2_decap_8 FILLER_41_341 ();
 sg13g2_decap_8 FILLER_41_348 ();
 sg13g2_decap_8 FILLER_41_355 ();
 sg13g2_decap_8 FILLER_41_362 ();
 sg13g2_decap_8 FILLER_41_369 ();
 sg13g2_decap_8 FILLER_41_376 ();
 sg13g2_decap_8 FILLER_41_383 ();
 sg13g2_decap_8 FILLER_41_390 ();
 sg13g2_decap_8 FILLER_41_397 ();
 sg13g2_decap_8 FILLER_41_404 ();
 sg13g2_decap_8 FILLER_41_411 ();
 sg13g2_decap_8 FILLER_41_418 ();
 sg13g2_decap_8 FILLER_41_425 ();
 sg13g2_decap_8 FILLER_41_432 ();
 sg13g2_decap_8 FILLER_41_439 ();
 sg13g2_decap_8 FILLER_41_446 ();
 sg13g2_decap_8 FILLER_41_453 ();
 sg13g2_decap_8 FILLER_41_460 ();
 sg13g2_decap_8 FILLER_41_467 ();
 sg13g2_decap_8 FILLER_41_474 ();
 sg13g2_decap_8 FILLER_41_481 ();
 sg13g2_decap_8 FILLER_41_488 ();
 sg13g2_decap_8 FILLER_41_495 ();
 sg13g2_decap_8 FILLER_41_502 ();
 sg13g2_decap_8 FILLER_41_509 ();
 sg13g2_decap_8 FILLER_41_516 ();
 sg13g2_decap_8 FILLER_41_523 ();
 sg13g2_decap_8 FILLER_41_530 ();
 sg13g2_decap_8 FILLER_41_537 ();
 sg13g2_decap_8 FILLER_41_544 ();
 sg13g2_decap_8 FILLER_41_551 ();
 sg13g2_decap_8 FILLER_41_558 ();
 sg13g2_decap_8 FILLER_41_565 ();
 sg13g2_decap_8 FILLER_41_572 ();
 sg13g2_decap_8 FILLER_41_579 ();
 sg13g2_decap_8 FILLER_41_586 ();
 sg13g2_decap_8 FILLER_41_593 ();
 sg13g2_decap_8 FILLER_41_600 ();
 sg13g2_decap_8 FILLER_41_607 ();
 sg13g2_decap_8 FILLER_41_614 ();
 sg13g2_decap_8 FILLER_41_621 ();
 sg13g2_decap_8 FILLER_41_628 ();
 sg13g2_decap_8 FILLER_41_635 ();
 sg13g2_decap_8 FILLER_41_642 ();
 sg13g2_decap_8 FILLER_41_649 ();
 sg13g2_decap_8 FILLER_41_656 ();
 sg13g2_decap_8 FILLER_41_663 ();
 sg13g2_decap_8 FILLER_41_670 ();
 sg13g2_decap_8 FILLER_41_677 ();
 sg13g2_decap_8 FILLER_41_684 ();
 sg13g2_decap_8 FILLER_41_691 ();
 sg13g2_decap_8 FILLER_41_698 ();
 sg13g2_decap_8 FILLER_41_705 ();
 sg13g2_decap_8 FILLER_41_712 ();
 sg13g2_decap_8 FILLER_41_719 ();
 sg13g2_decap_8 FILLER_41_726 ();
 sg13g2_decap_8 FILLER_41_733 ();
 sg13g2_decap_8 FILLER_41_740 ();
 sg13g2_decap_8 FILLER_41_747 ();
 sg13g2_decap_8 FILLER_41_754 ();
 sg13g2_decap_8 FILLER_41_761 ();
 sg13g2_decap_8 FILLER_41_768 ();
 sg13g2_decap_8 FILLER_41_775 ();
 sg13g2_decap_8 FILLER_41_782 ();
 sg13g2_decap_8 FILLER_41_789 ();
 sg13g2_decap_8 FILLER_41_796 ();
 sg13g2_decap_8 FILLER_41_803 ();
 sg13g2_decap_8 FILLER_41_810 ();
 sg13g2_decap_8 FILLER_41_817 ();
 sg13g2_decap_8 FILLER_41_824 ();
 sg13g2_decap_8 FILLER_41_831 ();
 sg13g2_decap_8 FILLER_41_838 ();
 sg13g2_decap_8 FILLER_41_845 ();
 sg13g2_decap_8 FILLER_41_852 ();
 sg13g2_decap_8 FILLER_41_859 ();
 sg13g2_decap_8 FILLER_41_866 ();
 sg13g2_decap_8 FILLER_41_873 ();
 sg13g2_decap_8 FILLER_41_880 ();
 sg13g2_decap_8 FILLER_41_887 ();
 sg13g2_decap_8 FILLER_41_894 ();
 sg13g2_decap_8 FILLER_41_901 ();
 sg13g2_decap_8 FILLER_41_908 ();
 sg13g2_decap_8 FILLER_41_915 ();
 sg13g2_decap_8 FILLER_41_922 ();
 sg13g2_decap_8 FILLER_41_929 ();
 sg13g2_decap_8 FILLER_41_936 ();
 sg13g2_decap_8 FILLER_41_943 ();
 sg13g2_decap_8 FILLER_41_950 ();
 sg13g2_decap_8 FILLER_41_957 ();
 sg13g2_decap_8 FILLER_41_964 ();
 sg13g2_decap_8 FILLER_41_971 ();
 sg13g2_decap_8 FILLER_41_978 ();
 sg13g2_decap_8 FILLER_41_985 ();
 sg13g2_decap_8 FILLER_41_992 ();
 sg13g2_decap_8 FILLER_41_999 ();
 sg13g2_decap_8 FILLER_41_1006 ();
 sg13g2_decap_8 FILLER_41_1013 ();
 sg13g2_decap_8 FILLER_41_1020 ();
 sg13g2_fill_2 FILLER_41_1027 ();
 sg13g2_decap_8 FILLER_42_5 ();
 sg13g2_decap_8 FILLER_42_12 ();
 sg13g2_decap_8 FILLER_42_19 ();
 sg13g2_decap_8 FILLER_42_26 ();
 sg13g2_decap_8 FILLER_42_33 ();
 sg13g2_decap_8 FILLER_42_40 ();
 sg13g2_decap_8 FILLER_42_47 ();
 sg13g2_decap_8 FILLER_42_54 ();
 sg13g2_decap_8 FILLER_42_61 ();
 sg13g2_decap_8 FILLER_42_68 ();
 sg13g2_decap_8 FILLER_42_75 ();
 sg13g2_decap_8 FILLER_42_82 ();
 sg13g2_decap_8 FILLER_42_89 ();
 sg13g2_decap_8 FILLER_42_96 ();
 sg13g2_decap_8 FILLER_42_103 ();
 sg13g2_decap_8 FILLER_42_110 ();
 sg13g2_decap_8 FILLER_42_117 ();
 sg13g2_decap_8 FILLER_42_124 ();
 sg13g2_decap_8 FILLER_42_131 ();
 sg13g2_decap_8 FILLER_42_138 ();
 sg13g2_decap_8 FILLER_42_145 ();
 sg13g2_decap_8 FILLER_42_152 ();
 sg13g2_decap_8 FILLER_42_159 ();
 sg13g2_decap_8 FILLER_42_166 ();
 sg13g2_decap_8 FILLER_42_173 ();
 sg13g2_decap_8 FILLER_42_180 ();
 sg13g2_decap_8 FILLER_42_187 ();
 sg13g2_decap_8 FILLER_42_194 ();
 sg13g2_decap_8 FILLER_42_201 ();
 sg13g2_decap_8 FILLER_42_208 ();
 sg13g2_decap_8 FILLER_42_215 ();
 sg13g2_decap_8 FILLER_42_222 ();
 sg13g2_decap_8 FILLER_42_229 ();
 sg13g2_decap_8 FILLER_42_236 ();
 sg13g2_decap_8 FILLER_42_243 ();
 sg13g2_decap_8 FILLER_42_250 ();
 sg13g2_decap_8 FILLER_42_257 ();
 sg13g2_decap_8 FILLER_42_264 ();
 sg13g2_decap_8 FILLER_42_271 ();
 sg13g2_decap_8 FILLER_42_278 ();
 sg13g2_decap_8 FILLER_42_285 ();
 sg13g2_decap_8 FILLER_42_292 ();
 sg13g2_decap_8 FILLER_42_299 ();
 sg13g2_decap_8 FILLER_42_306 ();
 sg13g2_decap_8 FILLER_42_313 ();
 sg13g2_decap_8 FILLER_42_320 ();
 sg13g2_decap_8 FILLER_42_327 ();
 sg13g2_decap_8 FILLER_42_334 ();
 sg13g2_decap_8 FILLER_42_341 ();
 sg13g2_decap_8 FILLER_42_348 ();
 sg13g2_decap_8 FILLER_42_355 ();
 sg13g2_decap_8 FILLER_42_362 ();
 sg13g2_decap_8 FILLER_42_369 ();
 sg13g2_decap_8 FILLER_42_376 ();
 sg13g2_decap_8 FILLER_42_383 ();
 sg13g2_decap_8 FILLER_42_390 ();
 sg13g2_decap_8 FILLER_42_397 ();
 sg13g2_decap_8 FILLER_42_404 ();
 sg13g2_decap_8 FILLER_42_411 ();
 sg13g2_decap_8 FILLER_42_418 ();
 sg13g2_decap_8 FILLER_42_425 ();
 sg13g2_decap_8 FILLER_42_432 ();
 sg13g2_decap_8 FILLER_42_439 ();
 sg13g2_decap_8 FILLER_42_446 ();
 sg13g2_decap_8 FILLER_42_453 ();
 sg13g2_decap_8 FILLER_42_460 ();
 sg13g2_decap_8 FILLER_42_467 ();
 sg13g2_decap_8 FILLER_42_474 ();
 sg13g2_decap_8 FILLER_42_481 ();
 sg13g2_decap_8 FILLER_42_488 ();
 sg13g2_decap_8 FILLER_42_495 ();
 sg13g2_decap_8 FILLER_42_502 ();
 sg13g2_decap_8 FILLER_42_509 ();
 sg13g2_decap_8 FILLER_42_516 ();
 sg13g2_decap_8 FILLER_42_523 ();
 sg13g2_decap_8 FILLER_42_530 ();
 sg13g2_decap_8 FILLER_42_537 ();
 sg13g2_decap_8 FILLER_42_544 ();
 sg13g2_decap_8 FILLER_42_551 ();
 sg13g2_decap_8 FILLER_42_558 ();
 sg13g2_decap_8 FILLER_42_565 ();
 sg13g2_decap_8 FILLER_42_572 ();
 sg13g2_decap_8 FILLER_42_579 ();
 sg13g2_decap_8 FILLER_42_586 ();
 sg13g2_decap_8 FILLER_42_593 ();
 sg13g2_decap_8 FILLER_42_600 ();
 sg13g2_decap_8 FILLER_42_607 ();
 sg13g2_decap_8 FILLER_42_614 ();
 sg13g2_decap_8 FILLER_42_621 ();
 sg13g2_decap_8 FILLER_42_628 ();
 sg13g2_decap_8 FILLER_42_635 ();
 sg13g2_decap_8 FILLER_42_642 ();
 sg13g2_decap_8 FILLER_42_649 ();
 sg13g2_decap_8 FILLER_42_656 ();
 sg13g2_decap_8 FILLER_42_663 ();
 sg13g2_decap_8 FILLER_42_670 ();
 sg13g2_decap_8 FILLER_42_677 ();
 sg13g2_decap_8 FILLER_42_684 ();
 sg13g2_decap_8 FILLER_42_691 ();
 sg13g2_decap_8 FILLER_42_698 ();
 sg13g2_decap_8 FILLER_42_705 ();
 sg13g2_decap_8 FILLER_42_712 ();
 sg13g2_decap_8 FILLER_42_719 ();
 sg13g2_decap_8 FILLER_42_726 ();
 sg13g2_decap_8 FILLER_42_733 ();
 sg13g2_decap_8 FILLER_42_740 ();
 sg13g2_decap_8 FILLER_42_747 ();
 sg13g2_decap_8 FILLER_42_754 ();
 sg13g2_decap_8 FILLER_42_761 ();
 sg13g2_decap_8 FILLER_42_768 ();
 sg13g2_decap_8 FILLER_42_775 ();
 sg13g2_decap_8 FILLER_42_782 ();
 sg13g2_decap_8 FILLER_42_789 ();
 sg13g2_decap_8 FILLER_42_796 ();
 sg13g2_decap_8 FILLER_42_803 ();
 sg13g2_decap_8 FILLER_42_810 ();
 sg13g2_decap_8 FILLER_42_817 ();
 sg13g2_decap_8 FILLER_42_824 ();
 sg13g2_decap_8 FILLER_42_831 ();
 sg13g2_decap_8 FILLER_42_838 ();
 sg13g2_decap_8 FILLER_42_845 ();
 sg13g2_decap_8 FILLER_42_852 ();
 sg13g2_decap_8 FILLER_42_859 ();
 sg13g2_decap_8 FILLER_42_866 ();
 sg13g2_decap_8 FILLER_42_873 ();
 sg13g2_decap_8 FILLER_42_880 ();
 sg13g2_decap_8 FILLER_42_887 ();
 sg13g2_decap_8 FILLER_42_894 ();
 sg13g2_decap_8 FILLER_42_901 ();
 sg13g2_decap_8 FILLER_42_908 ();
 sg13g2_decap_8 FILLER_42_915 ();
 sg13g2_decap_8 FILLER_42_922 ();
 sg13g2_decap_8 FILLER_42_929 ();
 sg13g2_decap_8 FILLER_42_936 ();
 sg13g2_decap_8 FILLER_42_943 ();
 sg13g2_decap_8 FILLER_42_950 ();
 sg13g2_decap_8 FILLER_42_957 ();
 sg13g2_decap_8 FILLER_42_964 ();
 sg13g2_decap_8 FILLER_42_971 ();
 sg13g2_decap_8 FILLER_42_978 ();
 sg13g2_decap_8 FILLER_42_985 ();
 sg13g2_decap_8 FILLER_42_992 ();
 sg13g2_decap_8 FILLER_42_999 ();
 sg13g2_decap_8 FILLER_42_1006 ();
 sg13g2_decap_8 FILLER_42_1013 ();
 sg13g2_decap_8 FILLER_42_1020 ();
 sg13g2_fill_2 FILLER_42_1027 ();
 sg13g2_decap_8 FILLER_43_5 ();
 sg13g2_decap_8 FILLER_43_12 ();
 sg13g2_decap_8 FILLER_43_19 ();
 sg13g2_decap_8 FILLER_43_26 ();
 sg13g2_decap_8 FILLER_43_33 ();
 sg13g2_decap_8 FILLER_43_40 ();
 sg13g2_decap_8 FILLER_43_47 ();
 sg13g2_decap_8 FILLER_43_54 ();
 sg13g2_decap_8 FILLER_43_61 ();
 sg13g2_decap_8 FILLER_43_68 ();
 sg13g2_decap_8 FILLER_43_75 ();
 sg13g2_decap_8 FILLER_43_82 ();
 sg13g2_decap_8 FILLER_43_89 ();
 sg13g2_decap_8 FILLER_43_96 ();
 sg13g2_decap_8 FILLER_43_103 ();
 sg13g2_decap_8 FILLER_43_110 ();
 sg13g2_decap_8 FILLER_43_117 ();
 sg13g2_decap_8 FILLER_43_124 ();
 sg13g2_decap_8 FILLER_43_131 ();
 sg13g2_decap_8 FILLER_43_138 ();
 sg13g2_decap_8 FILLER_43_145 ();
 sg13g2_decap_8 FILLER_43_152 ();
 sg13g2_decap_8 FILLER_43_159 ();
 sg13g2_decap_8 FILLER_43_166 ();
 sg13g2_decap_8 FILLER_43_173 ();
 sg13g2_decap_8 FILLER_43_180 ();
 sg13g2_decap_8 FILLER_43_187 ();
 sg13g2_decap_8 FILLER_43_194 ();
 sg13g2_decap_8 FILLER_43_201 ();
 sg13g2_decap_8 FILLER_43_208 ();
 sg13g2_decap_8 FILLER_43_215 ();
 sg13g2_decap_8 FILLER_43_222 ();
 sg13g2_decap_8 FILLER_43_229 ();
 sg13g2_decap_8 FILLER_43_236 ();
 sg13g2_decap_8 FILLER_43_243 ();
 sg13g2_decap_8 FILLER_43_250 ();
 sg13g2_decap_8 FILLER_43_257 ();
 sg13g2_decap_8 FILLER_43_264 ();
 sg13g2_decap_8 FILLER_43_271 ();
 sg13g2_decap_8 FILLER_43_278 ();
 sg13g2_decap_8 FILLER_43_285 ();
 sg13g2_decap_8 FILLER_43_292 ();
 sg13g2_decap_8 FILLER_43_299 ();
 sg13g2_decap_8 FILLER_43_306 ();
 sg13g2_decap_8 FILLER_43_313 ();
 sg13g2_decap_8 FILLER_43_320 ();
 sg13g2_decap_8 FILLER_43_327 ();
 sg13g2_decap_8 FILLER_43_334 ();
 sg13g2_decap_8 FILLER_43_341 ();
 sg13g2_decap_8 FILLER_43_348 ();
 sg13g2_decap_8 FILLER_43_355 ();
 sg13g2_decap_8 FILLER_43_362 ();
 sg13g2_decap_8 FILLER_43_369 ();
 sg13g2_decap_8 FILLER_43_376 ();
 sg13g2_decap_8 FILLER_43_383 ();
 sg13g2_decap_8 FILLER_43_390 ();
 sg13g2_decap_8 FILLER_43_397 ();
 sg13g2_decap_8 FILLER_43_404 ();
 sg13g2_decap_8 FILLER_43_411 ();
 sg13g2_decap_8 FILLER_43_418 ();
 sg13g2_decap_8 FILLER_43_425 ();
 sg13g2_decap_8 FILLER_43_432 ();
 sg13g2_decap_8 FILLER_43_439 ();
 sg13g2_decap_8 FILLER_43_446 ();
 sg13g2_decap_8 FILLER_43_453 ();
 sg13g2_decap_8 FILLER_43_460 ();
 sg13g2_decap_8 FILLER_43_467 ();
 sg13g2_decap_8 FILLER_43_474 ();
 sg13g2_decap_8 FILLER_43_481 ();
 sg13g2_decap_8 FILLER_43_488 ();
 sg13g2_decap_8 FILLER_43_495 ();
 sg13g2_decap_8 FILLER_43_502 ();
 sg13g2_decap_8 FILLER_43_509 ();
 sg13g2_decap_8 FILLER_43_516 ();
 sg13g2_decap_8 FILLER_43_523 ();
 sg13g2_decap_8 FILLER_43_530 ();
 sg13g2_decap_8 FILLER_43_537 ();
 sg13g2_decap_8 FILLER_43_544 ();
 sg13g2_decap_8 FILLER_43_551 ();
 sg13g2_decap_8 FILLER_43_558 ();
 sg13g2_decap_8 FILLER_43_565 ();
 sg13g2_decap_8 FILLER_43_572 ();
 sg13g2_decap_8 FILLER_43_579 ();
 sg13g2_decap_8 FILLER_43_586 ();
 sg13g2_decap_8 FILLER_43_593 ();
 sg13g2_decap_8 FILLER_43_600 ();
 sg13g2_decap_8 FILLER_43_607 ();
 sg13g2_decap_8 FILLER_43_614 ();
 sg13g2_decap_8 FILLER_43_621 ();
 sg13g2_decap_8 FILLER_43_628 ();
 sg13g2_decap_8 FILLER_43_635 ();
 sg13g2_decap_8 FILLER_43_642 ();
 sg13g2_decap_8 FILLER_43_649 ();
 sg13g2_decap_8 FILLER_43_656 ();
 sg13g2_decap_8 FILLER_43_663 ();
 sg13g2_decap_8 FILLER_43_670 ();
 sg13g2_decap_8 FILLER_43_677 ();
 sg13g2_decap_8 FILLER_43_684 ();
 sg13g2_decap_8 FILLER_43_691 ();
 sg13g2_decap_8 FILLER_43_698 ();
 sg13g2_decap_8 FILLER_43_705 ();
 sg13g2_decap_8 FILLER_43_712 ();
 sg13g2_decap_8 FILLER_43_719 ();
 sg13g2_decap_8 FILLER_43_726 ();
 sg13g2_decap_8 FILLER_43_733 ();
 sg13g2_decap_8 FILLER_43_740 ();
 sg13g2_decap_8 FILLER_43_747 ();
 sg13g2_decap_8 FILLER_43_754 ();
 sg13g2_decap_8 FILLER_43_761 ();
 sg13g2_decap_8 FILLER_43_768 ();
 sg13g2_decap_8 FILLER_43_775 ();
 sg13g2_decap_8 FILLER_43_782 ();
 sg13g2_decap_8 FILLER_43_789 ();
 sg13g2_decap_8 FILLER_43_796 ();
 sg13g2_decap_8 FILLER_43_803 ();
 sg13g2_decap_8 FILLER_43_810 ();
 sg13g2_decap_8 FILLER_43_817 ();
 sg13g2_decap_8 FILLER_43_824 ();
 sg13g2_decap_8 FILLER_43_831 ();
 sg13g2_decap_8 FILLER_43_838 ();
 sg13g2_decap_8 FILLER_43_845 ();
 sg13g2_decap_8 FILLER_43_852 ();
 sg13g2_decap_8 FILLER_43_859 ();
 sg13g2_decap_8 FILLER_43_866 ();
 sg13g2_decap_8 FILLER_43_873 ();
 sg13g2_decap_8 FILLER_43_880 ();
 sg13g2_decap_8 FILLER_43_887 ();
 sg13g2_decap_8 FILLER_43_894 ();
 sg13g2_decap_8 FILLER_43_901 ();
 sg13g2_decap_8 FILLER_43_908 ();
 sg13g2_decap_8 FILLER_43_915 ();
 sg13g2_decap_8 FILLER_43_922 ();
 sg13g2_decap_8 FILLER_43_929 ();
 sg13g2_decap_8 FILLER_43_936 ();
 sg13g2_decap_8 FILLER_43_943 ();
 sg13g2_decap_8 FILLER_43_950 ();
 sg13g2_decap_8 FILLER_43_957 ();
 sg13g2_decap_8 FILLER_43_964 ();
 sg13g2_decap_8 FILLER_43_971 ();
 sg13g2_decap_8 FILLER_43_978 ();
 sg13g2_decap_8 FILLER_43_985 ();
 sg13g2_decap_8 FILLER_43_992 ();
 sg13g2_decap_8 FILLER_43_999 ();
 sg13g2_decap_8 FILLER_43_1006 ();
 sg13g2_decap_8 FILLER_43_1013 ();
 sg13g2_decap_8 FILLER_43_1020 ();
 sg13g2_fill_2 FILLER_43_1027 ();
 sg13g2_decap_8 FILLER_44_5 ();
 sg13g2_decap_8 FILLER_44_12 ();
 sg13g2_decap_8 FILLER_44_19 ();
 sg13g2_decap_8 FILLER_44_26 ();
 sg13g2_decap_8 FILLER_44_33 ();
 sg13g2_decap_8 FILLER_44_40 ();
 sg13g2_decap_8 FILLER_44_47 ();
 sg13g2_decap_8 FILLER_44_54 ();
 sg13g2_decap_8 FILLER_44_61 ();
 sg13g2_decap_8 FILLER_44_68 ();
 sg13g2_decap_8 FILLER_44_75 ();
 sg13g2_decap_8 FILLER_44_82 ();
 sg13g2_decap_8 FILLER_44_89 ();
 sg13g2_decap_8 FILLER_44_96 ();
 sg13g2_decap_8 FILLER_44_103 ();
 sg13g2_decap_8 FILLER_44_110 ();
 sg13g2_decap_8 FILLER_44_117 ();
 sg13g2_decap_8 FILLER_44_124 ();
 sg13g2_decap_8 FILLER_44_131 ();
 sg13g2_decap_8 FILLER_44_138 ();
 sg13g2_decap_8 FILLER_44_145 ();
 sg13g2_decap_8 FILLER_44_152 ();
 sg13g2_decap_8 FILLER_44_159 ();
 sg13g2_decap_8 FILLER_44_166 ();
 sg13g2_decap_8 FILLER_44_173 ();
 sg13g2_decap_8 FILLER_44_180 ();
 sg13g2_decap_8 FILLER_44_187 ();
 sg13g2_decap_8 FILLER_44_194 ();
 sg13g2_decap_8 FILLER_44_201 ();
 sg13g2_decap_8 FILLER_44_208 ();
 sg13g2_decap_8 FILLER_44_215 ();
 sg13g2_decap_8 FILLER_44_222 ();
 sg13g2_decap_8 FILLER_44_229 ();
 sg13g2_decap_8 FILLER_44_236 ();
 sg13g2_decap_8 FILLER_44_243 ();
 sg13g2_decap_8 FILLER_44_250 ();
 sg13g2_decap_8 FILLER_44_257 ();
 sg13g2_decap_8 FILLER_44_264 ();
 sg13g2_decap_8 FILLER_44_271 ();
 sg13g2_decap_8 FILLER_44_278 ();
 sg13g2_decap_8 FILLER_44_285 ();
 sg13g2_decap_8 FILLER_44_292 ();
 sg13g2_decap_8 FILLER_44_299 ();
 sg13g2_decap_8 FILLER_44_306 ();
 sg13g2_decap_8 FILLER_44_313 ();
 sg13g2_decap_8 FILLER_44_320 ();
 sg13g2_decap_8 FILLER_44_327 ();
 sg13g2_decap_8 FILLER_44_334 ();
 sg13g2_decap_8 FILLER_44_341 ();
 sg13g2_decap_8 FILLER_44_348 ();
 sg13g2_decap_8 FILLER_44_355 ();
 sg13g2_decap_8 FILLER_44_362 ();
 sg13g2_decap_8 FILLER_44_369 ();
 sg13g2_decap_8 FILLER_44_376 ();
 sg13g2_decap_8 FILLER_44_383 ();
 sg13g2_decap_8 FILLER_44_390 ();
 sg13g2_decap_8 FILLER_44_397 ();
 sg13g2_decap_8 FILLER_44_404 ();
 sg13g2_decap_8 FILLER_44_411 ();
 sg13g2_decap_8 FILLER_44_418 ();
 sg13g2_decap_8 FILLER_44_425 ();
 sg13g2_decap_8 FILLER_44_432 ();
 sg13g2_decap_8 FILLER_44_439 ();
 sg13g2_decap_8 FILLER_44_446 ();
 sg13g2_decap_8 FILLER_44_453 ();
 sg13g2_decap_8 FILLER_44_460 ();
 sg13g2_decap_8 FILLER_44_467 ();
 sg13g2_decap_8 FILLER_44_474 ();
 sg13g2_decap_8 FILLER_44_481 ();
 sg13g2_decap_8 FILLER_44_488 ();
 sg13g2_decap_8 FILLER_44_495 ();
 sg13g2_decap_8 FILLER_44_502 ();
 sg13g2_decap_8 FILLER_44_509 ();
 sg13g2_decap_8 FILLER_44_516 ();
 sg13g2_decap_8 FILLER_44_523 ();
 sg13g2_decap_8 FILLER_44_530 ();
 sg13g2_decap_8 FILLER_44_537 ();
 sg13g2_decap_8 FILLER_44_544 ();
 sg13g2_decap_8 FILLER_44_551 ();
 sg13g2_decap_8 FILLER_44_558 ();
 sg13g2_decap_8 FILLER_44_565 ();
 sg13g2_decap_8 FILLER_44_572 ();
 sg13g2_decap_8 FILLER_44_579 ();
 sg13g2_decap_8 FILLER_44_586 ();
 sg13g2_decap_8 FILLER_44_593 ();
 sg13g2_decap_8 FILLER_44_600 ();
 sg13g2_decap_8 FILLER_44_607 ();
 sg13g2_decap_8 FILLER_44_614 ();
 sg13g2_decap_8 FILLER_44_621 ();
 sg13g2_decap_8 FILLER_44_628 ();
 sg13g2_decap_8 FILLER_44_635 ();
 sg13g2_decap_8 FILLER_44_642 ();
 sg13g2_decap_8 FILLER_44_649 ();
 sg13g2_decap_8 FILLER_44_656 ();
 sg13g2_decap_8 FILLER_44_663 ();
 sg13g2_decap_8 FILLER_44_670 ();
 sg13g2_decap_8 FILLER_44_677 ();
 sg13g2_decap_8 FILLER_44_684 ();
 sg13g2_decap_8 FILLER_44_691 ();
 sg13g2_decap_8 FILLER_44_698 ();
 sg13g2_decap_8 FILLER_44_705 ();
 sg13g2_decap_8 FILLER_44_712 ();
 sg13g2_decap_8 FILLER_44_719 ();
 sg13g2_decap_8 FILLER_44_726 ();
 sg13g2_decap_8 FILLER_44_733 ();
 sg13g2_decap_8 FILLER_44_740 ();
 sg13g2_decap_8 FILLER_44_747 ();
 sg13g2_decap_8 FILLER_44_754 ();
 sg13g2_decap_8 FILLER_44_761 ();
 sg13g2_decap_8 FILLER_44_768 ();
 sg13g2_decap_8 FILLER_44_775 ();
 sg13g2_decap_8 FILLER_44_782 ();
 sg13g2_decap_8 FILLER_44_789 ();
 sg13g2_decap_8 FILLER_44_796 ();
 sg13g2_decap_8 FILLER_44_803 ();
 sg13g2_decap_8 FILLER_44_810 ();
 sg13g2_decap_8 FILLER_44_817 ();
 sg13g2_decap_8 FILLER_44_824 ();
 sg13g2_decap_8 FILLER_44_831 ();
 sg13g2_decap_8 FILLER_44_838 ();
 sg13g2_decap_8 FILLER_44_845 ();
 sg13g2_decap_8 FILLER_44_852 ();
 sg13g2_decap_8 FILLER_44_859 ();
 sg13g2_decap_8 FILLER_44_866 ();
 sg13g2_decap_8 FILLER_44_873 ();
 sg13g2_decap_8 FILLER_44_880 ();
 sg13g2_decap_8 FILLER_44_887 ();
 sg13g2_decap_8 FILLER_44_894 ();
 sg13g2_decap_8 FILLER_44_901 ();
 sg13g2_decap_8 FILLER_44_908 ();
 sg13g2_decap_8 FILLER_44_915 ();
 sg13g2_decap_8 FILLER_44_922 ();
 sg13g2_decap_8 FILLER_44_929 ();
 sg13g2_decap_8 FILLER_44_936 ();
 sg13g2_decap_8 FILLER_44_943 ();
 sg13g2_decap_8 FILLER_44_950 ();
 sg13g2_decap_8 FILLER_44_957 ();
 sg13g2_decap_8 FILLER_44_964 ();
 sg13g2_decap_8 FILLER_44_971 ();
 sg13g2_decap_8 FILLER_44_978 ();
 sg13g2_decap_8 FILLER_44_985 ();
 sg13g2_decap_8 FILLER_44_992 ();
 sg13g2_decap_8 FILLER_44_999 ();
 sg13g2_decap_8 FILLER_44_1006 ();
 sg13g2_decap_8 FILLER_44_1013 ();
 sg13g2_decap_8 FILLER_44_1020 ();
 sg13g2_fill_2 FILLER_44_1027 ();
 sg13g2_decap_8 FILLER_45_5 ();
 sg13g2_decap_8 FILLER_45_12 ();
 sg13g2_decap_8 FILLER_45_19 ();
 sg13g2_decap_8 FILLER_45_26 ();
 sg13g2_decap_8 FILLER_45_33 ();
 sg13g2_decap_8 FILLER_45_40 ();
 sg13g2_decap_8 FILLER_45_47 ();
 sg13g2_decap_8 FILLER_45_54 ();
 sg13g2_decap_8 FILLER_45_61 ();
 sg13g2_decap_8 FILLER_45_68 ();
 sg13g2_decap_8 FILLER_45_75 ();
 sg13g2_decap_8 FILLER_45_82 ();
 sg13g2_decap_8 FILLER_45_89 ();
 sg13g2_decap_8 FILLER_45_96 ();
 sg13g2_decap_8 FILLER_45_103 ();
 sg13g2_decap_8 FILLER_45_110 ();
 sg13g2_decap_8 FILLER_45_117 ();
 sg13g2_decap_8 FILLER_45_124 ();
 sg13g2_decap_8 FILLER_45_131 ();
 sg13g2_decap_8 FILLER_45_138 ();
 sg13g2_decap_8 FILLER_45_145 ();
 sg13g2_decap_8 FILLER_45_152 ();
 sg13g2_decap_8 FILLER_45_159 ();
 sg13g2_decap_8 FILLER_45_166 ();
 sg13g2_decap_8 FILLER_45_173 ();
 sg13g2_decap_8 FILLER_45_180 ();
 sg13g2_decap_8 FILLER_45_187 ();
 sg13g2_decap_8 FILLER_45_194 ();
 sg13g2_decap_8 FILLER_45_201 ();
 sg13g2_decap_8 FILLER_45_208 ();
 sg13g2_decap_8 FILLER_45_215 ();
 sg13g2_decap_8 FILLER_45_222 ();
 sg13g2_decap_8 FILLER_45_229 ();
 sg13g2_decap_8 FILLER_45_236 ();
 sg13g2_decap_8 FILLER_45_243 ();
 sg13g2_decap_8 FILLER_45_250 ();
 sg13g2_decap_8 FILLER_45_257 ();
 sg13g2_decap_8 FILLER_45_264 ();
 sg13g2_decap_8 FILLER_45_271 ();
 sg13g2_decap_8 FILLER_45_278 ();
 sg13g2_decap_8 FILLER_45_285 ();
 sg13g2_decap_8 FILLER_45_292 ();
 sg13g2_decap_8 FILLER_45_299 ();
 sg13g2_decap_8 FILLER_45_306 ();
 sg13g2_decap_8 FILLER_45_313 ();
 sg13g2_decap_8 FILLER_45_320 ();
 sg13g2_decap_8 FILLER_45_327 ();
 sg13g2_decap_8 FILLER_45_334 ();
 sg13g2_decap_8 FILLER_45_341 ();
 sg13g2_decap_8 FILLER_45_348 ();
 sg13g2_decap_8 FILLER_45_355 ();
 sg13g2_decap_8 FILLER_45_362 ();
 sg13g2_decap_8 FILLER_45_369 ();
 sg13g2_decap_8 FILLER_45_376 ();
 sg13g2_decap_8 FILLER_45_383 ();
 sg13g2_decap_8 FILLER_45_390 ();
 sg13g2_decap_8 FILLER_45_397 ();
 sg13g2_decap_8 FILLER_45_404 ();
 sg13g2_decap_8 FILLER_45_411 ();
 sg13g2_decap_8 FILLER_45_418 ();
 sg13g2_decap_8 FILLER_45_425 ();
 sg13g2_decap_8 FILLER_45_432 ();
 sg13g2_decap_8 FILLER_45_439 ();
 sg13g2_decap_8 FILLER_45_446 ();
 sg13g2_decap_8 FILLER_45_453 ();
 sg13g2_decap_8 FILLER_45_460 ();
 sg13g2_decap_8 FILLER_45_467 ();
 sg13g2_decap_8 FILLER_45_474 ();
 sg13g2_decap_8 FILLER_45_481 ();
 sg13g2_decap_8 FILLER_45_488 ();
 sg13g2_decap_8 FILLER_45_495 ();
 sg13g2_decap_8 FILLER_45_502 ();
 sg13g2_decap_8 FILLER_45_509 ();
 sg13g2_decap_8 FILLER_45_516 ();
 sg13g2_decap_8 FILLER_45_523 ();
 sg13g2_decap_8 FILLER_45_530 ();
 sg13g2_decap_8 FILLER_45_537 ();
 sg13g2_decap_8 FILLER_45_544 ();
 sg13g2_decap_8 FILLER_45_551 ();
 sg13g2_decap_8 FILLER_45_558 ();
 sg13g2_decap_8 FILLER_45_565 ();
 sg13g2_decap_8 FILLER_45_572 ();
 sg13g2_decap_8 FILLER_45_579 ();
 sg13g2_decap_8 FILLER_45_586 ();
 sg13g2_decap_8 FILLER_45_593 ();
 sg13g2_decap_8 FILLER_45_600 ();
 sg13g2_decap_8 FILLER_45_607 ();
 sg13g2_decap_8 FILLER_45_614 ();
 sg13g2_decap_8 FILLER_45_621 ();
 sg13g2_decap_8 FILLER_45_628 ();
 sg13g2_decap_8 FILLER_45_635 ();
 sg13g2_decap_8 FILLER_45_642 ();
 sg13g2_decap_8 FILLER_45_649 ();
 sg13g2_decap_8 FILLER_45_656 ();
 sg13g2_decap_8 FILLER_45_663 ();
 sg13g2_decap_8 FILLER_45_670 ();
 sg13g2_decap_8 FILLER_45_677 ();
 sg13g2_decap_8 FILLER_45_684 ();
 sg13g2_decap_8 FILLER_45_691 ();
 sg13g2_decap_8 FILLER_45_698 ();
 sg13g2_decap_8 FILLER_45_705 ();
 sg13g2_decap_8 FILLER_45_712 ();
 sg13g2_decap_8 FILLER_45_719 ();
 sg13g2_decap_8 FILLER_45_726 ();
 sg13g2_decap_8 FILLER_45_733 ();
 sg13g2_decap_8 FILLER_45_740 ();
 sg13g2_decap_8 FILLER_45_747 ();
 sg13g2_decap_8 FILLER_45_754 ();
 sg13g2_decap_8 FILLER_45_761 ();
 sg13g2_decap_8 FILLER_45_768 ();
 sg13g2_decap_8 FILLER_45_775 ();
 sg13g2_decap_8 FILLER_45_782 ();
 sg13g2_decap_8 FILLER_45_789 ();
 sg13g2_decap_8 FILLER_45_796 ();
 sg13g2_decap_8 FILLER_45_803 ();
 sg13g2_decap_8 FILLER_45_810 ();
 sg13g2_decap_8 FILLER_45_817 ();
 sg13g2_decap_8 FILLER_45_824 ();
 sg13g2_decap_8 FILLER_45_831 ();
 sg13g2_decap_8 FILLER_45_838 ();
 sg13g2_decap_8 FILLER_45_845 ();
 sg13g2_decap_8 FILLER_45_852 ();
 sg13g2_decap_8 FILLER_45_859 ();
 sg13g2_decap_8 FILLER_45_866 ();
 sg13g2_decap_8 FILLER_45_873 ();
 sg13g2_decap_8 FILLER_45_880 ();
 sg13g2_decap_8 FILLER_45_887 ();
 sg13g2_decap_8 FILLER_45_894 ();
 sg13g2_decap_8 FILLER_45_901 ();
 sg13g2_decap_8 FILLER_45_908 ();
 sg13g2_decap_8 FILLER_45_915 ();
 sg13g2_decap_8 FILLER_45_922 ();
 sg13g2_decap_8 FILLER_45_929 ();
 sg13g2_decap_8 FILLER_45_936 ();
 sg13g2_decap_8 FILLER_45_943 ();
 sg13g2_decap_8 FILLER_45_950 ();
 sg13g2_decap_8 FILLER_45_957 ();
 sg13g2_decap_8 FILLER_45_964 ();
 sg13g2_decap_8 FILLER_45_971 ();
 sg13g2_decap_8 FILLER_45_978 ();
 sg13g2_decap_8 FILLER_45_985 ();
 sg13g2_decap_8 FILLER_45_992 ();
 sg13g2_decap_8 FILLER_45_999 ();
 sg13g2_decap_8 FILLER_45_1006 ();
 sg13g2_decap_8 FILLER_45_1013 ();
 sg13g2_decap_8 FILLER_45_1020 ();
 sg13g2_fill_2 FILLER_45_1027 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_28 ();
 sg13g2_decap_8 FILLER_46_35 ();
 sg13g2_decap_8 FILLER_46_42 ();
 sg13g2_decap_8 FILLER_46_49 ();
 sg13g2_decap_8 FILLER_46_56 ();
 sg13g2_decap_8 FILLER_46_63 ();
 sg13g2_decap_8 FILLER_46_70 ();
 sg13g2_decap_8 FILLER_46_77 ();
 sg13g2_decap_8 FILLER_46_84 ();
 sg13g2_decap_8 FILLER_46_91 ();
 sg13g2_decap_8 FILLER_46_98 ();
 sg13g2_decap_8 FILLER_46_105 ();
 sg13g2_decap_8 FILLER_46_112 ();
 sg13g2_decap_8 FILLER_46_119 ();
 sg13g2_decap_8 FILLER_46_126 ();
 sg13g2_decap_8 FILLER_46_133 ();
 sg13g2_decap_8 FILLER_46_140 ();
 sg13g2_decap_8 FILLER_46_147 ();
 sg13g2_decap_8 FILLER_46_154 ();
 sg13g2_decap_8 FILLER_46_161 ();
 sg13g2_decap_8 FILLER_46_168 ();
 sg13g2_decap_8 FILLER_46_175 ();
 sg13g2_decap_8 FILLER_46_182 ();
 sg13g2_decap_8 FILLER_46_189 ();
 sg13g2_decap_8 FILLER_46_196 ();
 sg13g2_decap_8 FILLER_46_203 ();
 sg13g2_decap_8 FILLER_46_210 ();
 sg13g2_decap_8 FILLER_46_217 ();
 sg13g2_decap_8 FILLER_46_224 ();
 sg13g2_decap_8 FILLER_46_231 ();
 sg13g2_decap_8 FILLER_46_238 ();
 sg13g2_decap_8 FILLER_46_245 ();
 sg13g2_decap_8 FILLER_46_252 ();
 sg13g2_decap_8 FILLER_46_259 ();
 sg13g2_decap_8 FILLER_46_266 ();
 sg13g2_decap_8 FILLER_46_273 ();
 sg13g2_decap_8 FILLER_46_280 ();
 sg13g2_decap_8 FILLER_46_287 ();
 sg13g2_decap_8 FILLER_46_294 ();
 sg13g2_decap_8 FILLER_46_301 ();
 sg13g2_decap_8 FILLER_46_308 ();
 sg13g2_decap_8 FILLER_46_315 ();
 sg13g2_decap_8 FILLER_46_322 ();
 sg13g2_decap_8 FILLER_46_329 ();
 sg13g2_decap_8 FILLER_46_336 ();
 sg13g2_decap_8 FILLER_46_343 ();
 sg13g2_decap_8 FILLER_46_350 ();
 sg13g2_decap_8 FILLER_46_357 ();
 sg13g2_decap_8 FILLER_46_364 ();
 sg13g2_decap_8 FILLER_46_371 ();
 sg13g2_decap_8 FILLER_46_378 ();
 sg13g2_decap_8 FILLER_46_385 ();
 sg13g2_decap_8 FILLER_46_392 ();
 sg13g2_decap_8 FILLER_46_399 ();
 sg13g2_decap_8 FILLER_46_406 ();
 sg13g2_decap_8 FILLER_46_413 ();
 sg13g2_decap_8 FILLER_46_420 ();
 sg13g2_decap_8 FILLER_46_427 ();
 sg13g2_decap_8 FILLER_46_434 ();
 sg13g2_decap_8 FILLER_46_441 ();
 sg13g2_decap_8 FILLER_46_448 ();
 sg13g2_decap_8 FILLER_46_455 ();
 sg13g2_decap_8 FILLER_46_462 ();
 sg13g2_decap_8 FILLER_46_469 ();
 sg13g2_decap_8 FILLER_46_476 ();
 sg13g2_decap_8 FILLER_46_483 ();
 sg13g2_decap_8 FILLER_46_490 ();
 sg13g2_decap_8 FILLER_46_497 ();
 sg13g2_decap_8 FILLER_46_504 ();
 sg13g2_decap_8 FILLER_46_511 ();
 sg13g2_decap_8 FILLER_46_518 ();
 sg13g2_decap_8 FILLER_46_525 ();
 sg13g2_decap_8 FILLER_46_532 ();
 sg13g2_decap_8 FILLER_46_539 ();
 sg13g2_decap_8 FILLER_46_546 ();
 sg13g2_decap_8 FILLER_46_553 ();
 sg13g2_decap_8 FILLER_46_560 ();
 sg13g2_decap_8 FILLER_46_567 ();
 sg13g2_decap_8 FILLER_46_574 ();
 sg13g2_decap_8 FILLER_46_581 ();
 sg13g2_decap_8 FILLER_46_588 ();
 sg13g2_decap_8 FILLER_46_595 ();
 sg13g2_decap_8 FILLER_46_602 ();
 sg13g2_decap_8 FILLER_46_609 ();
 sg13g2_decap_8 FILLER_46_616 ();
 sg13g2_decap_8 FILLER_46_623 ();
 sg13g2_decap_8 FILLER_46_630 ();
 sg13g2_decap_8 FILLER_46_637 ();
 sg13g2_decap_8 FILLER_46_644 ();
 sg13g2_decap_8 FILLER_46_651 ();
 sg13g2_decap_8 FILLER_46_658 ();
 sg13g2_decap_8 FILLER_46_665 ();
 sg13g2_decap_8 FILLER_46_672 ();
 sg13g2_decap_8 FILLER_46_679 ();
 sg13g2_decap_8 FILLER_46_686 ();
 sg13g2_decap_8 FILLER_46_693 ();
 sg13g2_decap_8 FILLER_46_700 ();
 sg13g2_decap_8 FILLER_46_707 ();
 sg13g2_decap_8 FILLER_46_714 ();
 sg13g2_decap_8 FILLER_46_721 ();
 sg13g2_decap_8 FILLER_46_728 ();
 sg13g2_decap_8 FILLER_46_735 ();
 sg13g2_decap_8 FILLER_46_742 ();
 sg13g2_decap_8 FILLER_46_749 ();
 sg13g2_decap_8 FILLER_46_756 ();
 sg13g2_decap_8 FILLER_46_763 ();
 sg13g2_decap_8 FILLER_46_770 ();
 sg13g2_decap_8 FILLER_46_777 ();
 sg13g2_decap_8 FILLER_46_784 ();
 sg13g2_decap_8 FILLER_46_791 ();
 sg13g2_decap_8 FILLER_46_798 ();
 sg13g2_decap_8 FILLER_46_805 ();
 sg13g2_decap_8 FILLER_46_812 ();
 sg13g2_decap_8 FILLER_46_819 ();
 sg13g2_decap_8 FILLER_46_826 ();
 sg13g2_decap_8 FILLER_46_833 ();
 sg13g2_decap_8 FILLER_46_840 ();
 sg13g2_decap_8 FILLER_46_847 ();
 sg13g2_decap_8 FILLER_46_854 ();
 sg13g2_decap_8 FILLER_46_861 ();
 sg13g2_decap_8 FILLER_46_868 ();
 sg13g2_decap_8 FILLER_46_875 ();
 sg13g2_decap_8 FILLER_46_882 ();
 sg13g2_decap_8 FILLER_46_889 ();
 sg13g2_decap_8 FILLER_46_896 ();
 sg13g2_decap_8 FILLER_46_903 ();
 sg13g2_decap_8 FILLER_46_910 ();
 sg13g2_decap_8 FILLER_46_917 ();
 sg13g2_decap_8 FILLER_46_924 ();
 sg13g2_decap_8 FILLER_46_931 ();
 sg13g2_decap_8 FILLER_46_938 ();
 sg13g2_decap_8 FILLER_46_945 ();
 sg13g2_decap_8 FILLER_46_952 ();
 sg13g2_decap_8 FILLER_46_959 ();
 sg13g2_decap_8 FILLER_46_966 ();
 sg13g2_decap_8 FILLER_46_973 ();
 sg13g2_decap_8 FILLER_46_980 ();
 sg13g2_decap_8 FILLER_46_987 ();
 sg13g2_decap_8 FILLER_46_994 ();
 sg13g2_decap_8 FILLER_46_1001 ();
 sg13g2_decap_8 FILLER_46_1008 ();
 sg13g2_decap_8 FILLER_46_1015 ();
 sg13g2_decap_8 FILLER_46_1022 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_8 FILLER_47_35 ();
 sg13g2_decap_8 FILLER_47_42 ();
 sg13g2_decap_8 FILLER_47_49 ();
 sg13g2_decap_8 FILLER_47_56 ();
 sg13g2_decap_8 FILLER_47_63 ();
 sg13g2_decap_8 FILLER_47_70 ();
 sg13g2_decap_8 FILLER_47_77 ();
 sg13g2_decap_8 FILLER_47_84 ();
 sg13g2_decap_8 FILLER_47_91 ();
 sg13g2_decap_8 FILLER_47_98 ();
 sg13g2_decap_8 FILLER_47_105 ();
 sg13g2_decap_8 FILLER_47_112 ();
 sg13g2_decap_8 FILLER_47_119 ();
 sg13g2_decap_8 FILLER_47_126 ();
 sg13g2_decap_8 FILLER_47_133 ();
 sg13g2_decap_8 FILLER_47_140 ();
 sg13g2_decap_8 FILLER_47_147 ();
 sg13g2_decap_8 FILLER_47_154 ();
 sg13g2_decap_8 FILLER_47_161 ();
 sg13g2_decap_8 FILLER_47_168 ();
 sg13g2_decap_8 FILLER_47_175 ();
 sg13g2_decap_8 FILLER_47_182 ();
 sg13g2_decap_8 FILLER_47_189 ();
 sg13g2_decap_8 FILLER_47_196 ();
 sg13g2_decap_8 FILLER_47_203 ();
 sg13g2_decap_8 FILLER_47_210 ();
 sg13g2_decap_8 FILLER_47_217 ();
 sg13g2_decap_8 FILLER_47_224 ();
 sg13g2_decap_8 FILLER_47_231 ();
 sg13g2_decap_8 FILLER_47_238 ();
 sg13g2_decap_8 FILLER_47_245 ();
 sg13g2_decap_8 FILLER_47_252 ();
 sg13g2_decap_8 FILLER_47_259 ();
 sg13g2_decap_8 FILLER_47_266 ();
 sg13g2_decap_8 FILLER_47_273 ();
 sg13g2_decap_8 FILLER_47_280 ();
 sg13g2_decap_8 FILLER_47_287 ();
 sg13g2_decap_8 FILLER_47_294 ();
 sg13g2_decap_8 FILLER_47_301 ();
 sg13g2_decap_8 FILLER_47_308 ();
 sg13g2_decap_8 FILLER_47_315 ();
 sg13g2_decap_8 FILLER_47_322 ();
 sg13g2_decap_8 FILLER_47_329 ();
 sg13g2_decap_8 FILLER_47_336 ();
 sg13g2_decap_8 FILLER_47_343 ();
 sg13g2_decap_8 FILLER_47_350 ();
 sg13g2_decap_8 FILLER_47_357 ();
 sg13g2_decap_8 FILLER_47_364 ();
 sg13g2_decap_8 FILLER_47_371 ();
 sg13g2_decap_8 FILLER_47_378 ();
 sg13g2_decap_8 FILLER_47_385 ();
 sg13g2_decap_8 FILLER_47_392 ();
 sg13g2_decap_8 FILLER_47_399 ();
 sg13g2_decap_8 FILLER_47_406 ();
 sg13g2_decap_8 FILLER_47_413 ();
 sg13g2_decap_8 FILLER_47_420 ();
 sg13g2_decap_8 FILLER_47_427 ();
 sg13g2_decap_8 FILLER_47_434 ();
 sg13g2_decap_8 FILLER_47_441 ();
 sg13g2_decap_8 FILLER_47_448 ();
 sg13g2_decap_8 FILLER_47_455 ();
 sg13g2_decap_8 FILLER_47_462 ();
 sg13g2_decap_8 FILLER_47_469 ();
 sg13g2_decap_8 FILLER_47_476 ();
 sg13g2_decap_8 FILLER_47_483 ();
 sg13g2_decap_8 FILLER_47_490 ();
 sg13g2_decap_8 FILLER_47_497 ();
 sg13g2_decap_8 FILLER_47_504 ();
 sg13g2_decap_8 FILLER_47_511 ();
 sg13g2_decap_8 FILLER_47_518 ();
 sg13g2_decap_8 FILLER_47_525 ();
 sg13g2_decap_8 FILLER_47_532 ();
 sg13g2_decap_8 FILLER_47_539 ();
 sg13g2_decap_8 FILLER_47_546 ();
 sg13g2_decap_8 FILLER_47_553 ();
 sg13g2_decap_8 FILLER_47_560 ();
 sg13g2_decap_8 FILLER_47_567 ();
 sg13g2_decap_8 FILLER_47_574 ();
 sg13g2_decap_8 FILLER_47_581 ();
 sg13g2_decap_8 FILLER_47_588 ();
 sg13g2_decap_8 FILLER_47_595 ();
 sg13g2_decap_8 FILLER_47_602 ();
 sg13g2_decap_8 FILLER_47_609 ();
 sg13g2_decap_8 FILLER_47_616 ();
 sg13g2_decap_8 FILLER_47_623 ();
 sg13g2_decap_8 FILLER_47_630 ();
 sg13g2_decap_8 FILLER_47_637 ();
 sg13g2_decap_8 FILLER_47_644 ();
 sg13g2_decap_8 FILLER_47_651 ();
 sg13g2_decap_8 FILLER_47_658 ();
 sg13g2_decap_8 FILLER_47_665 ();
 sg13g2_decap_8 FILLER_47_672 ();
 sg13g2_decap_8 FILLER_47_679 ();
 sg13g2_decap_8 FILLER_47_686 ();
 sg13g2_decap_8 FILLER_47_693 ();
 sg13g2_decap_8 FILLER_47_700 ();
 sg13g2_decap_8 FILLER_47_707 ();
 sg13g2_decap_8 FILLER_47_714 ();
 sg13g2_decap_8 FILLER_47_721 ();
 sg13g2_decap_8 FILLER_47_728 ();
 sg13g2_decap_8 FILLER_47_735 ();
 sg13g2_decap_8 FILLER_47_742 ();
 sg13g2_decap_8 FILLER_47_749 ();
 sg13g2_decap_8 FILLER_47_756 ();
 sg13g2_decap_8 FILLER_47_763 ();
 sg13g2_decap_8 FILLER_47_770 ();
 sg13g2_decap_8 FILLER_47_777 ();
 sg13g2_decap_8 FILLER_47_784 ();
 sg13g2_decap_8 FILLER_47_791 ();
 sg13g2_decap_8 FILLER_47_798 ();
 sg13g2_decap_8 FILLER_47_805 ();
 sg13g2_decap_8 FILLER_47_812 ();
 sg13g2_decap_8 FILLER_47_819 ();
 sg13g2_decap_8 FILLER_47_826 ();
 sg13g2_decap_8 FILLER_47_833 ();
 sg13g2_decap_8 FILLER_47_840 ();
 sg13g2_decap_8 FILLER_47_847 ();
 sg13g2_decap_8 FILLER_47_854 ();
 sg13g2_decap_8 FILLER_47_861 ();
 sg13g2_decap_8 FILLER_47_868 ();
 sg13g2_decap_8 FILLER_47_875 ();
 sg13g2_decap_8 FILLER_47_882 ();
 sg13g2_decap_8 FILLER_47_889 ();
 sg13g2_decap_8 FILLER_47_896 ();
 sg13g2_decap_8 FILLER_47_903 ();
 sg13g2_decap_8 FILLER_47_910 ();
 sg13g2_decap_8 FILLER_47_917 ();
 sg13g2_decap_8 FILLER_47_924 ();
 sg13g2_decap_8 FILLER_47_931 ();
 sg13g2_decap_8 FILLER_47_938 ();
 sg13g2_decap_8 FILLER_47_945 ();
 sg13g2_decap_8 FILLER_47_952 ();
 sg13g2_decap_8 FILLER_47_959 ();
 sg13g2_decap_8 FILLER_47_966 ();
 sg13g2_decap_8 FILLER_47_973 ();
 sg13g2_decap_8 FILLER_47_980 ();
 sg13g2_decap_8 FILLER_47_987 ();
 sg13g2_decap_8 FILLER_47_994 ();
 sg13g2_decap_8 FILLER_47_1001 ();
 sg13g2_decap_8 FILLER_47_1008 ();
 sg13g2_decap_8 FILLER_47_1015 ();
 sg13g2_decap_8 FILLER_47_1022 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_decap_8 FILLER_48_42 ();
 sg13g2_decap_8 FILLER_48_49 ();
 sg13g2_decap_8 FILLER_48_56 ();
 sg13g2_decap_8 FILLER_48_63 ();
 sg13g2_decap_8 FILLER_48_70 ();
 sg13g2_decap_8 FILLER_48_77 ();
 sg13g2_decap_8 FILLER_48_84 ();
 sg13g2_decap_8 FILLER_48_91 ();
 sg13g2_decap_8 FILLER_48_98 ();
 sg13g2_decap_8 FILLER_48_105 ();
 sg13g2_decap_8 FILLER_48_112 ();
 sg13g2_decap_8 FILLER_48_119 ();
 sg13g2_decap_8 FILLER_48_126 ();
 sg13g2_decap_8 FILLER_48_133 ();
 sg13g2_decap_8 FILLER_48_140 ();
 sg13g2_decap_8 FILLER_48_147 ();
 sg13g2_decap_8 FILLER_48_154 ();
 sg13g2_decap_8 FILLER_48_161 ();
 sg13g2_decap_8 FILLER_48_168 ();
 sg13g2_decap_8 FILLER_48_175 ();
 sg13g2_decap_8 FILLER_48_182 ();
 sg13g2_decap_8 FILLER_48_189 ();
 sg13g2_decap_8 FILLER_48_196 ();
 sg13g2_decap_8 FILLER_48_203 ();
 sg13g2_decap_8 FILLER_48_210 ();
 sg13g2_decap_8 FILLER_48_217 ();
 sg13g2_decap_8 FILLER_48_224 ();
 sg13g2_decap_8 FILLER_48_231 ();
 sg13g2_decap_8 FILLER_48_238 ();
 sg13g2_decap_8 FILLER_48_245 ();
 sg13g2_decap_8 FILLER_48_252 ();
 sg13g2_decap_8 FILLER_48_259 ();
 sg13g2_decap_8 FILLER_48_266 ();
 sg13g2_decap_8 FILLER_48_273 ();
 sg13g2_decap_8 FILLER_48_280 ();
 sg13g2_decap_8 FILLER_48_287 ();
 sg13g2_decap_8 FILLER_48_294 ();
 sg13g2_decap_8 FILLER_48_301 ();
 sg13g2_decap_8 FILLER_48_308 ();
 sg13g2_decap_8 FILLER_48_315 ();
 sg13g2_decap_8 FILLER_48_322 ();
 sg13g2_decap_8 FILLER_48_329 ();
 sg13g2_decap_8 FILLER_48_336 ();
 sg13g2_decap_8 FILLER_48_343 ();
 sg13g2_decap_8 FILLER_48_350 ();
 sg13g2_decap_8 FILLER_48_357 ();
 sg13g2_decap_8 FILLER_48_364 ();
 sg13g2_decap_8 FILLER_48_371 ();
 sg13g2_decap_8 FILLER_48_378 ();
 sg13g2_decap_8 FILLER_48_385 ();
 sg13g2_decap_8 FILLER_48_392 ();
 sg13g2_decap_8 FILLER_48_399 ();
 sg13g2_decap_8 FILLER_48_406 ();
 sg13g2_decap_8 FILLER_48_413 ();
 sg13g2_decap_8 FILLER_48_420 ();
 sg13g2_decap_8 FILLER_48_427 ();
 sg13g2_decap_8 FILLER_48_434 ();
 sg13g2_decap_8 FILLER_48_441 ();
 sg13g2_decap_8 FILLER_48_448 ();
 sg13g2_decap_8 FILLER_48_455 ();
 sg13g2_decap_8 FILLER_48_462 ();
 sg13g2_decap_8 FILLER_48_469 ();
 sg13g2_decap_8 FILLER_48_476 ();
 sg13g2_decap_8 FILLER_48_483 ();
 sg13g2_decap_8 FILLER_48_490 ();
 sg13g2_decap_8 FILLER_48_497 ();
 sg13g2_decap_8 FILLER_48_504 ();
 sg13g2_decap_8 FILLER_48_511 ();
 sg13g2_decap_8 FILLER_48_518 ();
 sg13g2_decap_8 FILLER_48_525 ();
 sg13g2_decap_8 FILLER_48_532 ();
 sg13g2_decap_8 FILLER_48_539 ();
 sg13g2_decap_8 FILLER_48_546 ();
 sg13g2_decap_8 FILLER_48_553 ();
 sg13g2_decap_8 FILLER_48_560 ();
 sg13g2_decap_8 FILLER_48_567 ();
 sg13g2_decap_8 FILLER_48_574 ();
 sg13g2_decap_8 FILLER_48_581 ();
 sg13g2_decap_8 FILLER_48_588 ();
 sg13g2_decap_8 FILLER_48_595 ();
 sg13g2_decap_8 FILLER_48_602 ();
 sg13g2_decap_8 FILLER_48_609 ();
 sg13g2_decap_8 FILLER_48_616 ();
 sg13g2_decap_8 FILLER_48_623 ();
 sg13g2_decap_8 FILLER_48_630 ();
 sg13g2_decap_8 FILLER_48_637 ();
 sg13g2_decap_8 FILLER_48_644 ();
 sg13g2_decap_8 FILLER_48_651 ();
 sg13g2_decap_8 FILLER_48_658 ();
 sg13g2_decap_8 FILLER_48_665 ();
 sg13g2_decap_8 FILLER_48_672 ();
 sg13g2_decap_8 FILLER_48_679 ();
 sg13g2_decap_8 FILLER_48_686 ();
 sg13g2_decap_8 FILLER_48_693 ();
 sg13g2_decap_8 FILLER_48_700 ();
 sg13g2_decap_8 FILLER_48_707 ();
 sg13g2_decap_8 FILLER_48_714 ();
 sg13g2_decap_8 FILLER_48_721 ();
 sg13g2_decap_8 FILLER_48_728 ();
 sg13g2_decap_8 FILLER_48_735 ();
 sg13g2_decap_8 FILLER_48_742 ();
 sg13g2_decap_8 FILLER_48_749 ();
 sg13g2_decap_8 FILLER_48_756 ();
 sg13g2_decap_8 FILLER_48_763 ();
 sg13g2_decap_8 FILLER_48_770 ();
 sg13g2_decap_8 FILLER_48_777 ();
 sg13g2_decap_8 FILLER_48_784 ();
 sg13g2_decap_8 FILLER_48_791 ();
 sg13g2_decap_8 FILLER_48_798 ();
 sg13g2_decap_8 FILLER_48_805 ();
 sg13g2_decap_8 FILLER_48_812 ();
 sg13g2_decap_8 FILLER_48_819 ();
 sg13g2_decap_8 FILLER_48_826 ();
 sg13g2_decap_8 FILLER_48_833 ();
 sg13g2_decap_8 FILLER_48_840 ();
 sg13g2_decap_8 FILLER_48_847 ();
 sg13g2_decap_8 FILLER_48_854 ();
 sg13g2_decap_8 FILLER_48_861 ();
 sg13g2_decap_8 FILLER_48_868 ();
 sg13g2_decap_8 FILLER_48_875 ();
 sg13g2_decap_8 FILLER_48_882 ();
 sg13g2_decap_8 FILLER_48_889 ();
 sg13g2_decap_8 FILLER_48_896 ();
 sg13g2_decap_8 FILLER_48_903 ();
 sg13g2_decap_8 FILLER_48_910 ();
 sg13g2_decap_8 FILLER_48_917 ();
 sg13g2_decap_8 FILLER_48_924 ();
 sg13g2_decap_8 FILLER_48_931 ();
 sg13g2_decap_8 FILLER_48_938 ();
 sg13g2_decap_8 FILLER_48_945 ();
 sg13g2_decap_8 FILLER_48_952 ();
 sg13g2_decap_8 FILLER_48_959 ();
 sg13g2_decap_8 FILLER_48_966 ();
 sg13g2_decap_8 FILLER_48_973 ();
 sg13g2_decap_8 FILLER_48_980 ();
 sg13g2_decap_8 FILLER_48_987 ();
 sg13g2_decap_8 FILLER_48_994 ();
 sg13g2_decap_8 FILLER_48_1001 ();
 sg13g2_decap_8 FILLER_48_1008 ();
 sg13g2_decap_8 FILLER_48_1015 ();
 sg13g2_decap_8 FILLER_48_1022 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_8 FILLER_49_28 ();
 sg13g2_decap_8 FILLER_49_35 ();
 sg13g2_decap_8 FILLER_49_42 ();
 sg13g2_decap_8 FILLER_49_49 ();
 sg13g2_decap_8 FILLER_49_56 ();
 sg13g2_decap_8 FILLER_49_63 ();
 sg13g2_decap_8 FILLER_49_70 ();
 sg13g2_decap_8 FILLER_49_77 ();
 sg13g2_decap_8 FILLER_49_84 ();
 sg13g2_decap_8 FILLER_49_91 ();
 sg13g2_decap_8 FILLER_49_98 ();
 sg13g2_decap_8 FILLER_49_105 ();
 sg13g2_decap_8 FILLER_49_112 ();
 sg13g2_decap_8 FILLER_49_119 ();
 sg13g2_decap_8 FILLER_49_126 ();
 sg13g2_decap_8 FILLER_49_133 ();
 sg13g2_decap_8 FILLER_49_140 ();
 sg13g2_decap_8 FILLER_49_147 ();
 sg13g2_decap_8 FILLER_49_154 ();
 sg13g2_decap_8 FILLER_49_161 ();
 sg13g2_decap_8 FILLER_49_168 ();
 sg13g2_decap_8 FILLER_49_175 ();
 sg13g2_decap_8 FILLER_49_182 ();
 sg13g2_decap_8 FILLER_49_189 ();
 sg13g2_decap_8 FILLER_49_196 ();
 sg13g2_decap_8 FILLER_49_203 ();
 sg13g2_decap_8 FILLER_49_210 ();
 sg13g2_decap_8 FILLER_49_217 ();
 sg13g2_decap_8 FILLER_49_224 ();
 sg13g2_decap_8 FILLER_49_231 ();
 sg13g2_decap_8 FILLER_49_238 ();
 sg13g2_decap_8 FILLER_49_245 ();
 sg13g2_decap_8 FILLER_49_252 ();
 sg13g2_decap_8 FILLER_49_259 ();
 sg13g2_decap_8 FILLER_49_266 ();
 sg13g2_decap_8 FILLER_49_273 ();
 sg13g2_decap_8 FILLER_49_280 ();
 sg13g2_decap_8 FILLER_49_287 ();
 sg13g2_decap_8 FILLER_49_294 ();
 sg13g2_decap_8 FILLER_49_301 ();
 sg13g2_decap_8 FILLER_49_308 ();
 sg13g2_decap_8 FILLER_49_315 ();
 sg13g2_decap_8 FILLER_49_322 ();
 sg13g2_decap_8 FILLER_49_329 ();
 sg13g2_decap_8 FILLER_49_336 ();
 sg13g2_decap_8 FILLER_49_343 ();
 sg13g2_decap_8 FILLER_49_350 ();
 sg13g2_decap_8 FILLER_49_357 ();
 sg13g2_decap_8 FILLER_49_364 ();
 sg13g2_decap_8 FILLER_49_371 ();
 sg13g2_decap_8 FILLER_49_378 ();
 sg13g2_decap_8 FILLER_49_385 ();
 sg13g2_decap_8 FILLER_49_392 ();
 sg13g2_decap_8 FILLER_49_399 ();
 sg13g2_decap_8 FILLER_49_406 ();
 sg13g2_decap_8 FILLER_49_413 ();
 sg13g2_decap_8 FILLER_49_420 ();
 sg13g2_decap_8 FILLER_49_427 ();
 sg13g2_decap_8 FILLER_49_434 ();
 sg13g2_decap_8 FILLER_49_441 ();
 sg13g2_decap_8 FILLER_49_448 ();
 sg13g2_decap_8 FILLER_49_455 ();
 sg13g2_decap_8 FILLER_49_462 ();
 sg13g2_decap_8 FILLER_49_469 ();
 sg13g2_decap_8 FILLER_49_476 ();
 sg13g2_decap_8 FILLER_49_483 ();
 sg13g2_decap_8 FILLER_49_490 ();
 sg13g2_decap_8 FILLER_49_497 ();
 sg13g2_decap_8 FILLER_49_504 ();
 sg13g2_decap_8 FILLER_49_511 ();
 sg13g2_decap_8 FILLER_49_518 ();
 sg13g2_decap_8 FILLER_49_525 ();
 sg13g2_decap_8 FILLER_49_532 ();
 sg13g2_decap_8 FILLER_49_539 ();
 sg13g2_decap_8 FILLER_49_546 ();
 sg13g2_decap_8 FILLER_49_553 ();
 sg13g2_decap_8 FILLER_49_560 ();
 sg13g2_decap_8 FILLER_49_567 ();
 sg13g2_decap_8 FILLER_49_574 ();
 sg13g2_decap_8 FILLER_49_581 ();
 sg13g2_decap_8 FILLER_49_588 ();
 sg13g2_decap_8 FILLER_49_595 ();
 sg13g2_decap_8 FILLER_49_602 ();
 sg13g2_decap_8 FILLER_49_609 ();
 sg13g2_decap_8 FILLER_49_616 ();
 sg13g2_decap_8 FILLER_49_623 ();
 sg13g2_decap_8 FILLER_49_630 ();
 sg13g2_decap_8 FILLER_49_637 ();
 sg13g2_decap_8 FILLER_49_644 ();
 sg13g2_decap_8 FILLER_49_651 ();
 sg13g2_decap_8 FILLER_49_658 ();
 sg13g2_decap_8 FILLER_49_665 ();
 sg13g2_decap_8 FILLER_49_672 ();
 sg13g2_decap_8 FILLER_49_679 ();
 sg13g2_decap_8 FILLER_49_686 ();
 sg13g2_decap_8 FILLER_49_693 ();
 sg13g2_decap_8 FILLER_49_700 ();
 sg13g2_decap_8 FILLER_49_707 ();
 sg13g2_decap_8 FILLER_49_714 ();
 sg13g2_decap_8 FILLER_49_721 ();
 sg13g2_decap_8 FILLER_49_728 ();
 sg13g2_decap_8 FILLER_49_735 ();
 sg13g2_decap_8 FILLER_49_742 ();
 sg13g2_decap_8 FILLER_49_749 ();
 sg13g2_decap_8 FILLER_49_756 ();
 sg13g2_decap_8 FILLER_49_763 ();
 sg13g2_decap_8 FILLER_49_770 ();
 sg13g2_decap_8 FILLER_49_777 ();
 sg13g2_decap_8 FILLER_49_784 ();
 sg13g2_decap_8 FILLER_49_791 ();
 sg13g2_decap_8 FILLER_49_798 ();
 sg13g2_decap_8 FILLER_49_805 ();
 sg13g2_decap_8 FILLER_49_812 ();
 sg13g2_decap_8 FILLER_49_819 ();
 sg13g2_decap_8 FILLER_49_826 ();
 sg13g2_decap_8 FILLER_49_833 ();
 sg13g2_decap_8 FILLER_49_840 ();
 sg13g2_decap_8 FILLER_49_847 ();
 sg13g2_decap_8 FILLER_49_854 ();
 sg13g2_decap_8 FILLER_49_861 ();
 sg13g2_decap_8 FILLER_49_868 ();
 sg13g2_decap_8 FILLER_49_875 ();
 sg13g2_decap_8 FILLER_49_882 ();
 sg13g2_decap_8 FILLER_49_889 ();
 sg13g2_decap_8 FILLER_49_896 ();
 sg13g2_decap_8 FILLER_49_903 ();
 sg13g2_decap_8 FILLER_49_910 ();
 sg13g2_decap_8 FILLER_49_917 ();
 sg13g2_decap_8 FILLER_49_924 ();
 sg13g2_decap_8 FILLER_49_931 ();
 sg13g2_decap_8 FILLER_49_938 ();
 sg13g2_decap_8 FILLER_49_945 ();
 sg13g2_decap_8 FILLER_49_952 ();
 sg13g2_decap_8 FILLER_49_959 ();
 sg13g2_decap_8 FILLER_49_966 ();
 sg13g2_decap_8 FILLER_49_973 ();
 sg13g2_decap_8 FILLER_49_980 ();
 sg13g2_decap_8 FILLER_49_987 ();
 sg13g2_decap_8 FILLER_49_994 ();
 sg13g2_decap_8 FILLER_49_1001 ();
 sg13g2_decap_8 FILLER_49_1008 ();
 sg13g2_decap_8 FILLER_49_1015 ();
 sg13g2_decap_8 FILLER_49_1022 ();
 assign uio_oe[0] = net38;
 assign uio_oe[1] = net39;
 assign uio_oe[2] = net40;
 assign uio_oe[3] = net41;
 assign uio_oe[4] = net42;
 assign uio_oe[5] = net43;
 assign uio_oe[6] = net44;
 assign uio_oe[7] = net45;
 assign uio_out[4] = net33;
 assign uio_out[5] = net34;
 assign uio_out[6] = net35;
 assign uio_out[7] = net36;
endmodule
