* NGSPICE file created from heichips25_template.ext - technology: ihp-sg13g2

* Black-box entry subcircuit for sg13g2_decap_8 abstract view
.subckt sg13g2_decap_8 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_2 abstract view
.subckt sg13g2_fill_2 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dfrbpq_1 abstract view
.subckt sg13g2_dfrbpq_1 RESET_B VSS VDD D Q CLK
.ends

* Black-box entry subcircuit for sg13g2_or2_1 abstract view
.subckt sg13g2_or2_1 VSS VDD X B A
.ends

* Black-box entry subcircuit for sg13g2_decap_4 abstract view
.subckt sg13g2_decap_4 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a22oi_1 abstract view
.subckt sg13g2_a22oi_1 Y B1 B2 A2 A1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_1 abstract view
.subckt sg13g2_fill_1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_1 abstract view
.subckt sg13g2_buf_1 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and2_1 abstract view
.subckt sg13g2_and2_1 A B X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2b_1 abstract view
.subckt sg13g2_nor2b_1 A B_N Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_tiehi abstract view
.subckt sg13g2_tiehi VDD VSS L_HI
.ends

* Black-box entry subcircuit for sg13g2_inv_1 abstract view
.subckt sg13g2_inv_1 VDD Y A VSS
.ends

* Black-box entry subcircuit for sg13g2_a21o_1 abstract view
.subckt sg13g2_a21o_1 A2 A1 B1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand3_1 abstract view
.subckt sg13g2_nand3_1 B C A Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_xor2_1 abstract view
.subckt sg13g2_xor2_1 B A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2b_1 abstract view
.subckt sg13g2_nand2b_1 Y B A_N VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_tielo abstract view
.subckt sg13g2_tielo VDD VSS L_LO
.ends

* Black-box entry subcircuit for sg13g2_buf_8 abstract view
.subckt sg13g2_buf_8 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2_1 abstract view
.subckt sg13g2_nor2_1 A B Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2_2 abstract view
.subckt sg13g2_nand2_2 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2_1 abstract view
.subckt sg13g2_nand2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2b_2 abstract view
.subckt sg13g2_nor2b_2 A B_N Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_2 abstract view
.subckt sg13g2_buf_2 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_2 abstract view
.subckt sg13g2_inv_2 Y A VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_4 abstract view
.subckt sg13g2_inv_4 A Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dfrbpq_2 abstract view
.subckt sg13g2_dfrbpq_2 RESET_B VSS VDD D Q CLK
.ends

* Black-box entry subcircuit for sg13g2_nor3_1 abstract view
.subckt sg13g2_nor3_1 A B C Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_mux2_1 abstract view
.subckt sg13g2_mux2_1 A0 A1 S X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_o21ai_1 abstract view
.subckt sg13g2_o21ai_1 B1 VDD Y VSS A1 A2
.ends

* Black-box entry subcircuit for sg13g2_dlygate4sd3_1 abstract view
.subckt sg13g2_dlygate4sd3_1 A VDD VSS X
.ends

* Black-box entry subcircuit for sg13g2_xnor2_1 abstract view
.subckt sg13g2_xnor2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand4_1 abstract view
.subckt sg13g2_nand4_1 B C A Y VDD VSS D
.ends

* Black-box entry subcircuit for sg13g2_nand3b_1 abstract view
.subckt sg13g2_nand3b_1 B C Y VDD VSS A_N
.ends

* Black-box entry subcircuit for sg13g2_nor2_2 abstract view
.subckt sg13g2_nor2_2 A B Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21oi_2 abstract view
.subckt sg13g2_a21oi_2 VSS VDD B1 Y A2 A1
.ends

* Black-box entry subcircuit for sg13g2_nor4_1 abstract view
.subckt sg13g2_nor4_1 A B C D Y VDD VSS
.ends

.subckt heichips25_template VGND VPWR clk ena rst_n ui_in[0] ui_in[1] ui_in[2] ui_in[3]
+ ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4]
+ uio_in[5] uio_in[6] uio_in[7] uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4]
+ uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4]
+ uio_out[5] uio_out[6] uio_out[7] uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4]
+ uo_out[5] uo_out[6] uo_out[7]
XFILLER_27_406 VPWR VGND sg13g2_decap_8
XFILLER_28_918 VPWR VGND sg13g2_decap_8
XFILLER_36_19 VPWR VGND sg13g2_decap_8
XFILLER_35_472 VPWR VGND sg13g2_decap_8
XFILLER_36_984 VPWR VGND sg13g2_decap_8
XFILLER_23_634 VPWR VGND sg13g2_decap_8
XFILLER_22_144 VPWR VGND sg13g2_decap_8
XFILLER_22_166 VPWR VGND sg13g2_decap_8
XFILLER_7_7 VPWR VGND sg13g2_decap_8
XFILLER_18_417 VPWR VGND sg13g2_decap_8
XFILLER_45_236 VPWR VGND sg13g2_decap_8
XFILLER_27_973 VPWR VGND sg13g2_decap_8
XFILLER_14_612 VPWR VGND sg13g2_decap_8
XFILLER_26_74 VPWR VGND sg13g2_decap_8
XFILLER_26_483 VPWR VGND sg13g2_decap_8
XFILLER_42_943 VPWR VGND sg13g2_decap_8
XFILLER_41_453 VPWR VGND sg13g2_decap_8
XFILLER_13_144 VPWR VGND sg13g2_decap_8
XFILLER_14_689 VPWR VGND sg13g2_decap_8
XFILLER_42_40 VPWR VGND sg13g2_decap_8
XFILLER_9_137 VPWR VGND sg13g2_decap_8
XFILLER_10_851 VPWR VGND sg13g2_decap_8
XFILLER_6_844 VPWR VGND sg13g2_decap_8
XFILLER_5_354 VPWR VGND sg13g2_decap_8
XFILLER_1_560 VPWR VGND sg13g2_decap_8
XFILLER_3_67 VPWR VGND sg13g2_decap_8
XFILLER_49_553 VPWR VGND sg13g2_decap_8
XFILLER_37_748 VPWR VGND sg13g2_decap_8
XFILLER_36_247 VPWR VGND sg13g2_decap_8
XFILLER_17_483 VPWR VGND sg13g2_decap_8
XFILLER_18_984 VPWR VGND sg13g2_decap_8
XFILLER_33_943 VPWR VGND sg13g2_decap_8
XFILLER_32_453 VPWR VGND sg13g2_decap_8
XFILLER_41_1013 VPWR VGND sg13g2_decap_8
XFILLER_28_715 VPWR VGND sg13g2_decap_8
XFILLER_27_203 VPWR VGND sg13g2_decap_8
XFILLER_24_921 VPWR VGND sg13g2_decap_8
XFILLER_36_781 VPWR VGND sg13g2_decap_8
XFILLER_23_431 VPWR VGND sg13g2_decap_8
XFILLER_24_998 VPWR VGND sg13g2_decap_8
XFILLER_11_648 VPWR VGND sg13g2_decap_8
XFILLER_10_158 VPWR VGND sg13g2_decap_8
XFILLER_12_32 VPWR VGND sg13g2_decap_8
XFILLER_5_4 VPWR VGND sg13g2_decap_8
XFILLER_3_858 VPWR VGND sg13g2_decap_8
XFILLER_2_368 VPWR VGND sg13g2_decap_8
XFILLER_18_214 VPWR VGND sg13g2_decap_8
XFILLER_19_748 VPWR VGND sg13g2_decap_8
XFILLER_46_567 VPWR VGND sg13g2_decap_8
XFILLER_37_84 VPWR VGND sg13g2_decap_8
XFILLER_15_910 VPWR VGND sg13g2_decap_8
XFILLER_27_770 VPWR VGND sg13g2_decap_8
XFILLER_42_740 VPWR VGND sg13g2_decap_8
XFILLER_15_987 VPWR VGND sg13g2_decap_8
XFILLER_18_1026 VPWR VGND sg13g2_fill_2
XFILLER_14_486 VPWR VGND sg13g2_decap_8
XFILLER_30_968 VPWR VGND sg13g2_decap_8
XFILLER_6_641 VPWR VGND sg13g2_decap_8
XFILLER_5_151 VPWR VGND sg13g2_decap_8
XFILLER_45_5 VPWR VGND sg13g2_decap_8
XFILLER_38_4 VPWR VGND sg13g2_decap_8
XFILLER_49_350 VPWR VGND sg13g2_decap_8
XFILLER_37_545 VPWR VGND sg13g2_decap_8
XFILLER_18_781 VPWR VGND sg13g2_decap_8
XFILLER_17_280 VPWR VGND sg13g2_decap_8
XFILLER_33_740 VPWR VGND sg13g2_decap_8
XFILLER_21_913 VPWR VGND sg13g2_decap_8
XFILLER_32_250 VPWR VGND sg13g2_decap_8
XFILLER_20_467 VPWR VGND sg13g2_decap_8
XFILLER_28_512 VPWR VGND sg13g2_decap_8
XFILLER_28_589 VPWR VGND sg13g2_decap_8
XFILLER_43_537 VPWR VGND sg13g2_decap_8
XFILLER_12_935 VPWR VGND sg13g2_decap_8
XFILLER_24_795 VPWR VGND sg13g2_decap_8
XFILLER_8_928 VPWR VGND sg13g2_decap_8
XFILLER_11_445 VPWR VGND sg13g2_decap_8
XFILLER_23_53 VPWR VGND sg13g2_decap_8
X_131_ net14 VGND VPWR mod1.qam16_mod.i_level\[2\] mod1.i_out_qam16\[2\] clknet_2_1__leaf_clk
+ sg13g2_dfrbpq_1
XFILLER_7_427 VPWR VGND sg13g2_decap_8
X_062_ VGND VPWR _037_ net10 net16 sg13g2_or2_1
XFILLER_48_1008 VPWR VGND sg13g2_decap_8
XFILLER_3_655 VPWR VGND sg13g2_decap_8
XFILLER_2_165 VPWR VGND sg13g2_decap_8
XFILLER_47_854 VPWR VGND sg13g2_decap_8
XFILLER_0_35 VPWR VGND sg13g2_decap_8
XFILLER_19_545 VPWR VGND sg13g2_decap_8
XFILLER_46_364 VPWR VGND sg13g2_decap_8
XFILLER_34_559 VPWR VGND sg13g2_decap_8
XFILLER_9_11 VPWR VGND sg13g2_decap_8
XFILLER_14_283 VPWR VGND sg13g2_decap_8
XFILLER_15_784 VPWR VGND sg13g2_decap_8
XFILLER_9_88 VPWR VGND sg13g2_decap_8
XFILLER_30_765 VPWR VGND sg13g2_decap_8
XFILLER_31_1023 VPWR VGND sg13g2_decap_4
XFILLER_7_994 VPWR VGND sg13g2_decap_8
XFILLER_29_0 VPWR VGND sg13g2_decap_8
XFILLER_37_342 VPWR VGND sg13g2_decap_8
XFILLER_38_876 VPWR VGND sg13g2_decap_8
XFILLER_44_19 VPWR VGND sg13g2_decap_8
XFILLER_25_537 VPWR VGND sg13g2_decap_8
XFILLER_21_710 VPWR VGND sg13g2_decap_8
XFILLER_20_242 VPWR VGND sg13g2_decap_8
XFILLER_21_787 VPWR VGND sg13g2_decap_8
XFILLER_0_658 VPWR VGND sg13g2_decap_8
XFILLER_18_53 VPWR VGND sg13g2_decap_8
XFILLER_28_342 VPWR VGND sg13g2_decap_4
XFILLER_29_865 VPWR VGND sg13g2_decap_8
XFILLER_44_824 VPWR VGND sg13g2_decap_8
XFILLER_28_375 VPWR VGND sg13g2_decap_8
XFILLER_43_334 VPWR VGND sg13g2_decap_8
XFILLER_16_559 VPWR VGND sg13g2_decap_8
XFILLER_12_732 VPWR VGND sg13g2_decap_8
XFILLER_24_592 VPWR VGND sg13g2_decap_8
XFILLER_34_96 VPWR VGND sg13g2_decap_8
XFILLER_8_725 VPWR VGND sg13g2_decap_8
XFILLER_11_242 VPWR VGND sg13g2_decap_8
XFILLER_7_224 VPWR VGND sg13g2_decap_8
X_114_ _004_ _027_ _028_ _025_ _023_ VPWR VGND sg13g2_a22oi_1
XFILLER_4_942 VPWR VGND sg13g2_decap_8
XFILLER_3_452 VPWR VGND sg13g2_decap_8
XFILLER_47_651 VPWR VGND sg13g2_decap_8
XFILLER_19_353 VPWR VGND sg13g2_decap_8
XFILLER_46_161 VPWR VGND sg13g2_decap_8
XFILLER_35_857 VPWR VGND sg13g2_decap_8
XFILLER_34_345 VPWR VGND sg13g2_decap_8
XFILLER_34_356 VPWR VGND sg13g2_fill_1
XFILLER_15_581 VPWR VGND sg13g2_decap_8
XFILLER_30_562 VPWR VGND sg13g2_decap_8
XFILLER_7_791 VPWR VGND sg13g2_decap_8
XFILLER_38_673 VPWR VGND sg13g2_decap_8
XFILLER_25_367 VPWR VGND sg13g2_decap_8
XFILLER_26_868 VPWR VGND sg13g2_decap_8
XFILLER_37_194 VPWR VGND sg13g2_decap_8
XFILLER_41_838 VPWR VGND sg13g2_decap_8
XFILLER_13_529 VPWR VGND sg13g2_decap_8
XFILLER_40_348 VPWR VGND sg13g2_decap_8
XFILLER_21_584 VPWR VGND sg13g2_decap_8
XFILLER_5_739 VPWR VGND sg13g2_decap_8
XFILLER_4_249 VPWR VGND sg13g2_decap_8
XFILLER_20_32 VPWR VGND sg13g2_decap_8
XFILLER_1_945 VPWR VGND sg13g2_decap_8
XFILLER_0_455 VPWR VGND sg13g2_decap_8
XFILLER_49_938 VPWR VGND sg13g2_decap_8
XFILLER_48_448 VPWR VGND sg13g2_decap_8
XFILLER_21_1011 VPWR VGND sg13g2_decap_8
XFILLER_29_63 VPWR VGND sg13g2_decap_8
XFILLER_29_662 VPWR VGND sg13g2_decap_8
XFILLER_45_40 VPWR VGND sg13g2_decap_8
XFILLER_44_621 VPWR VGND sg13g2_decap_8
XFILLER_16_312 VPWR VGND sg13g2_decap_8
XFILLER_28_183 VPWR VGND sg13g2_decap_8
XFILLER_43_131 VPWR VGND sg13g2_decap_8
XFILLER_16_356 VPWR VGND sg13g2_decap_8
XFILLER_17_868 VPWR VGND sg13g2_decap_8
XFILLER_44_698 VPWR VGND sg13g2_decap_8
XFILLER_32_838 VPWR VGND sg13g2_decap_8
XFILLER_31_337 VPWR VGND sg13g2_decap_8
XFILLER_8_522 VPWR VGND sg13g2_decap_8
XFILLER_8_599 VPWR VGND sg13g2_decap_8
XFILLER_6_67 VPWR VGND sg13g2_decap_8
XFILLER_6_1005 VPWR VGND sg13g2_decap_8
XFILLER_20_4 VPWR VGND sg13g2_decap_8
XFILLER_39_459 VPWR VGND sg13g2_decap_8
XFILLER_26_109 VPWR VGND sg13g2_decap_8
XFILLER_34_131 VPWR VGND sg13g2_decap_8
XFILLER_35_654 VPWR VGND sg13g2_decap_8
XFILLER_23_816 VPWR VGND sg13g2_decap_8
XFILLER_22_348 VPWR VGND sg13g2_decap_8
XFILLER_45_418 VPWR VGND sg13g2_decap_8
XFILLER_38_470 VPWR VGND sg13g2_decap_8
XFILLER_26_665 VPWR VGND sg13g2_decap_8
XFILLER_15_32 VPWR VGND sg13g2_decap_8
XFILLER_25_175 VPWR VGND sg13g2_decap_8
XFILLER_41_635 VPWR VGND sg13g2_decap_8
XFILLER_13_326 VPWR VGND sg13g2_decap_8
XFILLER_40_123 VPWR VGND sg13g2_decap_8
XFILLER_9_319 VPWR VGND sg13g2_decap_8
XFILLER_21_381 VPWR VGND sg13g2_decap_8
XFILLER_5_536 VPWR VGND sg13g2_decap_8
XFILLER_31_75 VPWR VGND sg13g2_decap_8
Xoutput20 net25 uo_out[0] VPWR VGND sg13g2_buf_1
XFILLER_1_742 VPWR VGND sg13g2_decap_8
XFILLER_0_252 VPWR VGND sg13g2_decap_8
XFILLER_49_735 VPWR VGND sg13g2_decap_8
XFILLER_48_245 VPWR VGND sg13g2_decap_8
XFILLER_17_665 VPWR VGND sg13g2_decap_8
XFILLER_45_985 VPWR VGND sg13g2_decap_8
XFILLER_44_495 VPWR VGND sg13g2_decap_8
XFILLER_16_186 VPWR VGND sg13g2_decap_8
XFILLER_32_635 VPWR VGND sg13g2_decap_8
XFILLER_31_145 VPWR VGND sg13g2_decap_8
XFILLER_13_893 VPWR VGND sg13g2_decap_8
XFILLER_9_886 VPWR VGND sg13g2_decap_8
XFILLER_8_396 VPWR VGND sg13g2_decap_8
XFILLER_39_256 VPWR VGND sg13g2_decap_8
XFILLER_36_963 VPWR VGND sg13g2_decap_8
XFILLER_23_613 VPWR VGND sg13g2_decap_8
XFILLER_35_451 VPWR VGND sg13g2_decap_8
XFILLER_22_123 VPWR VGND sg13g2_decap_8
XFILLER_46_749 VPWR VGND sg13g2_decap_8
XFILLER_45_215 VPWR VGND sg13g2_decap_8
XFILLER_27_952 VPWR VGND sg13g2_decap_8
XFILLER_42_922 VPWR VGND sg13g2_decap_8
XFILLER_26_53 VPWR VGND sg13g2_decap_8
XFILLER_26_462 VPWR VGND sg13g2_decap_8
XFILLER_41_432 VPWR VGND sg13g2_decap_8
XFILLER_13_123 VPWR VGND sg13g2_decap_8
XFILLER_42_999 VPWR VGND sg13g2_decap_8
XFILLER_9_116 VPWR VGND sg13g2_decap_8
XFILLER_14_668 VPWR VGND sg13g2_decap_8
XFILLER_10_830 VPWR VGND sg13g2_decap_8
XFILLER_42_96 VPWR VGND sg13g2_decap_8
XFILLER_6_823 VPWR VGND sg13g2_decap_8
XFILLER_5_333 VPWR VGND sg13g2_decap_8
XFILLER_3_46 VPWR VGND sg13g2_decap_8
XFILLER_49_532 VPWR VGND sg13g2_decap_8
XFILLER_3_1019 VPWR VGND sg13g2_decap_8
XFILLER_36_215 VPWR VGND sg13g2_decap_8
XFILLER_37_727 VPWR VGND sg13g2_decap_8
XFILLER_18_963 VPWR VGND sg13g2_decap_8
XFILLER_45_782 VPWR VGND sg13g2_decap_8
XFILLER_17_462 VPWR VGND sg13g2_decap_8
XFILLER_33_922 VPWR VGND sg13g2_decap_8
XFILLER_44_292 VPWR VGND sg13g2_decap_8
XFILLER_32_432 VPWR VGND sg13g2_decap_8
XFILLER_33_999 VPWR VGND sg13g2_decap_8
XFILLER_20_649 VPWR VGND sg13g2_decap_8
XFILLER_34_1021 VPWR VGND sg13g2_decap_8
XFILLER_13_690 VPWR VGND sg13g2_decap_8
XFILLER_9_683 VPWR VGND sg13g2_decap_8
XFILLER_8_193 VPWR VGND sg13g2_decap_8
XFILLER_27_259 VPWR VGND sg13g2_decap_8
XFILLER_43_719 VPWR VGND sg13g2_decap_8
XFILLER_24_900 VPWR VGND sg13g2_decap_8
XFILLER_36_760 VPWR VGND sg13g2_decap_8
XFILLER_42_229 VPWR VGND sg13g2_decap_8
XFILLER_23_410 VPWR VGND sg13g2_decap_8
XFILLER_35_292 VPWR VGND sg13g2_decap_4
XFILLER_24_977 VPWR VGND sg13g2_decap_8
XFILLER_11_627 VPWR VGND sg13g2_decap_8
XFILLER_23_487 VPWR VGND sg13g2_decap_8
XFILLER_10_137 VPWR VGND sg13g2_decap_8
XFILLER_7_609 VPWR VGND sg13g2_decap_8
XFILLER_12_11 VPWR VGND sg13g2_decap_8
XFILLER_12_88 VPWR VGND sg13g2_decap_8
XFILLER_3_837 VPWR VGND sg13g2_decap_8
XFILLER_2_347 VPWR VGND sg13g2_decap_8
XFILLER_19_727 VPWR VGND sg13g2_decap_8
XFILLER_46_546 VPWR VGND sg13g2_decap_8
XFILLER_37_63 VPWR VGND sg13g2_decap_8
XFILLER_26_281 VPWR VGND sg13g2_decap_8
XFILLER_33_229 VPWR VGND sg13g2_decap_8
XFILLER_14_465 VPWR VGND sg13g2_decap_8
XFILLER_15_966 VPWR VGND sg13g2_decap_8
XFILLER_18_1005 VPWR VGND sg13g2_decap_8
XFILLER_42_796 VPWR VGND sg13g2_decap_8
XFILLER_30_947 VPWR VGND sg13g2_decap_8
XFILLER_6_620 VPWR VGND sg13g2_decap_8
XFILLER_5_130 VPWR VGND sg13g2_decap_8
XFILLER_6_697 VPWR VGND sg13g2_decap_8
XFILLER_37_524 VPWR VGND sg13g2_decap_8
XFILLER_18_760 VPWR VGND sg13g2_decap_8
XFILLER_25_719 VPWR VGND sg13g2_decap_8
XFILLER_24_229 VPWR VGND sg13g2_decap_8
XFILLER_33_796 VPWR VGND sg13g2_decap_8
XFILLER_20_446 VPWR VGND sg13g2_decap_8
XFILLER_21_969 VPWR VGND sg13g2_decap_8
XFILLER_9_480 VPWR VGND sg13g2_decap_8
XFILLER_43_516 VPWR VGND sg13g2_decap_8
XFILLER_28_568 VPWR VGND sg13g2_decap_8
XFILLER_12_914 VPWR VGND sg13g2_decap_8
XFILLER_11_424 VPWR VGND sg13g2_decap_8
XFILLER_23_251 VPWR VGND sg13g2_decap_8
XFILLER_24_774 VPWR VGND sg13g2_decap_8
XFILLER_8_907 VPWR VGND sg13g2_decap_8
XFILLER_7_406 VPWR VGND sg13g2_decap_8
XFILLER_23_32 VPWR VGND sg13g2_decap_8
X_130_ net15 VGND VPWR _008_ mod1.i_out_8psk\[2\] clknet_2_3__leaf_clk sg13g2_dfrbpq_1
X_061_ net7 net6 _036_ VPWR VGND sg13g2_and2_1
XFILLER_3_634 VPWR VGND sg13g2_decap_8
XFILLER_2_144 VPWR VGND sg13g2_decap_8
XFILLER_47_833 VPWR VGND sg13g2_decap_8
XFILLER_48_84 VPWR VGND sg13g2_decap_8
XFILLER_19_524 VPWR VGND sg13g2_decap_8
XFILLER_46_343 VPWR VGND sg13g2_decap_8
XFILLER_0_14 VPWR VGND sg13g2_decap_8
XFILLER_34_538 VPWR VGND sg13g2_decap_8
XFILLER_15_763 VPWR VGND sg13g2_decap_8
XFILLER_14_262 VPWR VGND sg13g2_decap_8
XFILLER_42_593 VPWR VGND sg13g2_decap_8
XFILLER_9_67 VPWR VGND sg13g2_decap_8
XFILLER_30_744 VPWR VGND sg13g2_decap_8
XFILLER_31_1002 VPWR VGND sg13g2_decap_8
XFILLER_11_991 VPWR VGND sg13g2_decap_8
XFILLER_7_973 VPWR VGND sg13g2_decap_8
XFILLER_6_494 VPWR VGND sg13g2_decap_8
XFILLER_37_321 VPWR VGND sg13g2_decap_8
XFILLER_38_855 VPWR VGND sg13g2_decap_8
XFILLER_25_516 VPWR VGND sg13g2_decap_8
XFILLER_37_398 VPWR VGND sg13g2_decap_8
XFILLER_20_221 VPWR VGND sg13g2_decap_8
XFILLER_33_593 VPWR VGND sg13g2_decap_8
XFILLER_21_766 VPWR VGND sg13g2_decap_8
XFILLER_20_298 VPWR VGND sg13g2_decap_8
XFILLER_0_637 VPWR VGND sg13g2_decap_8
XFILLER_18_32 VPWR VGND sg13g2_decap_8
XFILLER_28_321 VPWR VGND sg13g2_decap_8
XFILLER_29_844 VPWR VGND sg13g2_decap_8
XFILLER_44_803 VPWR VGND sg13g2_decap_8
XFILLER_43_313 VPWR VGND sg13g2_decap_8
XFILLER_16_538 VPWR VGND sg13g2_decap_8
XFILLER_12_711 VPWR VGND sg13g2_decap_8
XFILLER_24_571 VPWR VGND sg13g2_decap_8
XFILLER_31_519 VPWR VGND sg13g2_decap_8
XFILLER_8_704 VPWR VGND sg13g2_decap_8
XFILLER_11_221 VPWR VGND sg13g2_decap_8
XFILLER_15_1008 VPWR VGND sg13g2_decap_8
XFILLER_34_75 VPWR VGND sg13g2_decap_8
XFILLER_7_203 VPWR VGND sg13g2_decap_8
XFILLER_12_788 VPWR VGND sg13g2_decap_8
XFILLER_11_298 VPWR VGND sg13g2_decap_8
X_113_ net20 net12 _028_ VPWR VGND sg13g2_nor2b_1
XFILLER_4_921 VPWR VGND sg13g2_decap_8
XFILLER_3_431 VPWR VGND sg13g2_decap_8
XFILLER_4_998 VPWR VGND sg13g2_decap_8
XFILLER_47_630 VPWR VGND sg13g2_decap_8
XFILLER_19_332 VPWR VGND sg13g2_decap_8
XFILLER_46_140 VPWR VGND sg13g2_decap_8
XFILLER_34_324 VPWR VGND sg13g2_decap_8
XFILLER_35_836 VPWR VGND sg13g2_decap_8
XFILLER_43_880 VPWR VGND sg13g2_decap_8
XFILLER_15_560 VPWR VGND sg13g2_decap_8
XFILLER_42_390 VPWR VGND sg13g2_decap_8
XFILLER_30_541 VPWR VGND sg13g2_decap_8
XFILLER_7_770 VPWR VGND sg13g2_decap_8
XFILLER_6_291 VPWR VGND sg13g2_decap_8
XFILLER_37_140 VPWR VGND sg13g2_decap_8
XFILLER_37_151 VPWR VGND sg13g2_fill_2
XFILLER_38_652 VPWR VGND sg13g2_decap_8
XFILLER_26_847 VPWR VGND sg13g2_decap_8
XFILLER_25_346 VPWR VGND sg13g2_decap_8
XFILLER_41_817 VPWR VGND sg13g2_decap_8
XFILLER_13_508 VPWR VGND sg13g2_decap_8
XFILLER_40_327 VPWR VGND sg13g2_decap_8
XFILLER_21_563 VPWR VGND sg13g2_decap_8
XFILLER_5_718 VPWR VGND sg13g2_decap_8
XFILLER_4_228 VPWR VGND sg13g2_decap_8
XFILLER_20_11 VPWR VGND sg13g2_decap_8
XFILLER_1_924 VPWR VGND sg13g2_decap_8
XFILLER_20_88 VPWR VGND sg13g2_decap_8
XFILLER_49_917 VPWR VGND sg13g2_decap_8
XFILLER_0_434 VPWR VGND sg13g2_decap_8
XFILLER_48_427 VPWR VGND sg13g2_decap_8
XFILLER_29_42 VPWR VGND sg13g2_decap_8
XFILLER_29_641 VPWR VGND sg13g2_decap_8
XFILLER_44_600 VPWR VGND sg13g2_decap_8
XFILLER_17_847 VPWR VGND sg13g2_decap_8
XFILLER_43_110 VPWR VGND sg13g2_decap_8
XFILLER_45_96 VPWR VGND sg13g2_decap_8
XFILLER_44_677 VPWR VGND sg13g2_decap_8
XFILLER_25_880 VPWR VGND sg13g2_decap_8
XFILLER_31_316 VPWR VGND sg13g2_decap_8
XFILLER_32_817 VPWR VGND sg13g2_decap_8
XFILLER_43_187 VPWR VGND sg13g2_decap_8
XFILLER_8_501 VPWR VGND sg13g2_decap_8
XFILLER_12_585 VPWR VGND sg13g2_decap_8
XFILLER_40_894 VPWR VGND sg13g2_decap_8
XFILLER_8_578 VPWR VGND sg13g2_decap_8
XFILLER_6_46 VPWR VGND sg13g2_decap_8
XFILLER_4_795 VPWR VGND sg13g2_decap_8
XFILLER_6_1028 VPWR VGND sg13g2_fill_1
XFILLER_13_4 VPWR VGND sg13g2_decap_8
XFILLER_39_438 VPWR VGND sg13g2_decap_8
XFILLER_48_994 VPWR VGND sg13g2_decap_8
XFILLER_19_151 VPWR VGND sg13g2_fill_2
XFILLER_35_633 VPWR VGND sg13g2_decap_8
XFILLER_34_110 VPWR VGND sg13g2_decap_8
XFILLER_22_327 VPWR VGND sg13g2_decap_8
XFILLER_34_187 VPWR VGND sg13g2_decap_8
XFILLER_34_198 VPWR VGND sg13g2_fill_2
XFILLER_31_883 VPWR VGND sg13g2_decap_8
Xheichips25_template_33 VPWR VGND uio_oe[0] sg13g2_tiehi
XFILLER_26_644 VPWR VGND sg13g2_decap_8
XFILLER_41_614 VPWR VGND sg13g2_decap_8
XFILLER_13_305 VPWR VGND sg13g2_decap_8
XFILLER_15_11 VPWR VGND sg13g2_decap_8
XFILLER_40_102 VPWR VGND sg13g2_decap_8
XFILLER_15_88 VPWR VGND sg13g2_decap_8
XFILLER_21_360 VPWR VGND sg13g2_decap_8
XFILLER_40_179 VPWR VGND sg13g2_decap_8
XFILLER_5_515 VPWR VGND sg13g2_decap_8
XFILLER_31_54 VPWR VGND sg13g2_decap_8
Xoutput21 net26 uo_out[1] VPWR VGND sg13g2_buf_1
XFILLER_1_721 VPWR VGND sg13g2_decap_8
XFILLER_49_714 VPWR VGND sg13g2_decap_8
XFILLER_0_231 VPWR VGND sg13g2_decap_8
XFILLER_48_224 VPWR VGND sg13g2_decap_8
XFILLER_1_798 VPWR VGND sg13g2_decap_8
XFILLER_37_909 VPWR VGND sg13g2_decap_8
XFILLER_45_964 VPWR VGND sg13g2_decap_8
XFILLER_17_644 VPWR VGND sg13g2_decap_8
XFILLER_44_474 VPWR VGND sg13g2_decap_8
XFILLER_16_165 VPWR VGND sg13g2_decap_8
XFILLER_32_614 VPWR VGND sg13g2_decap_8
XFILLER_31_124 VPWR VGND sg13g2_decap_8
XFILLER_13_872 VPWR VGND sg13g2_decap_8
XFILLER_12_382 VPWR VGND sg13g2_decap_8
XFILLER_9_865 VPWR VGND sg13g2_decap_8
XFILLER_40_691 VPWR VGND sg13g2_decap_8
XFILLER_8_375 VPWR VGND sg13g2_decap_8
XFILLER_4_592 VPWR VGND sg13g2_decap_8
XFILLER_39_235 VPWR VGND sg13g2_decap_8
XFILLER_48_791 VPWR VGND sg13g2_decap_8
XFILLER_35_430 VPWR VGND sg13g2_decap_8
XFILLER_36_942 VPWR VGND sg13g2_decap_8
XFILLER_22_102 VPWR VGND sg13g2_decap_8
XFILLER_11_809 VPWR VGND sg13g2_decap_8
XFILLER_23_669 VPWR VGND sg13g2_decap_8
XFILLER_10_319 VPWR VGND sg13g2_decap_8
XFILLER_31_680 VPWR VGND sg13g2_decap_8
XFILLER_2_529 VPWR VGND sg13g2_decap_8
XFILLER_19_909 VPWR VGND sg13g2_decap_8
XFILLER_46_728 VPWR VGND sg13g2_decap_8
XFILLER_26_32 VPWR VGND sg13g2_decap_8
XFILLER_27_931 VPWR VGND sg13g2_decap_8
XFILLER_42_901 VPWR VGND sg13g2_decap_8
XFILLER_26_441 VPWR VGND sg13g2_decap_8
XFILLER_41_411 VPWR VGND sg13g2_decap_8
XFILLER_13_102 VPWR VGND sg13g2_decap_8
XFILLER_14_647 VPWR VGND sg13g2_decap_8
XFILLER_42_978 VPWR VGND sg13g2_decap_8
XFILLER_41_488 VPWR VGND sg13g2_decap_8
XFILLER_13_179 VPWR VGND sg13g2_decap_8
XFILLER_42_75 VPWR VGND sg13g2_decap_8
XFILLER_6_802 VPWR VGND sg13g2_decap_8
XFILLER_21_190 VPWR VGND sg13g2_decap_8
XFILLER_5_312 VPWR VGND sg13g2_decap_8
XFILLER_10_886 VPWR VGND sg13g2_decap_8
XFILLER_6_879 VPWR VGND sg13g2_decap_8
XFILLER_5_389 VPWR VGND sg13g2_decap_8
XFILLER_3_25 VPWR VGND sg13g2_decap_8
XFILLER_49_511 VPWR VGND sg13g2_decap_8
XFILLER_1_595 VPWR VGND sg13g2_decap_8
XFILLER_37_706 VPWR VGND sg13g2_decap_8
XFILLER_49_588 VPWR VGND sg13g2_decap_8
XFILLER_18_942 VPWR VGND sg13g2_decap_8
XFILLER_45_761 VPWR VGND sg13g2_decap_8
XFILLER_17_441 VPWR VGND sg13g2_decap_8
XFILLER_33_901 VPWR VGND sg13g2_decap_8
XFILLER_44_271 VPWR VGND sg13g2_decap_8
XFILLER_32_411 VPWR VGND sg13g2_decap_8
XFILLER_33_978 VPWR VGND sg13g2_decap_8
XFILLER_34_1000 VPWR VGND sg13g2_decap_8
XFILLER_20_628 VPWR VGND sg13g2_decap_8
XFILLER_32_488 VPWR VGND sg13g2_decap_8
XFILLER_9_662 VPWR VGND sg13g2_decap_8
XFILLER_8_172 VPWR VGND sg13g2_decap_8
XFILLER_27_238 VPWR VGND sg13g2_decap_8
XFILLER_42_208 VPWR VGND sg13g2_decap_8
XFILLER_24_956 VPWR VGND sg13g2_decap_8
XFILLER_11_606 VPWR VGND sg13g2_decap_8
XFILLER_23_466 VPWR VGND sg13g2_decap_8
XFILLER_10_116 VPWR VGND sg13g2_decap_8
XFILLER_6_109 VPWR VGND sg13g2_decap_8
XFILLER_12_67 VPWR VGND sg13g2_decap_8
XFILLER_3_816 VPWR VGND sg13g2_decap_8
XFILLER_2_326 VPWR VGND sg13g2_decap_8
XFILLER_19_706 VPWR VGND sg13g2_decap_8
XFILLER_46_525 VPWR VGND sg13g2_decap_8
XFILLER_37_42 VPWR VGND sg13g2_decap_8
XFILLER_15_945 VPWR VGND sg13g2_decap_8
XFILLER_26_260 VPWR VGND sg13g2_decap_8
XFILLER_14_444 VPWR VGND sg13g2_decap_8
XFILLER_18_1028 VPWR VGND sg13g2_fill_1
XFILLER_42_775 VPWR VGND sg13g2_decap_8
XFILLER_30_926 VPWR VGND sg13g2_decap_8
XFILLER_41_263 VPWR VGND sg13g2_decap_8
XFILLER_41_285 VPWR VGND sg13g2_decap_8
XFILLER_10_683 VPWR VGND sg13g2_decap_8
XFILLER_6_676 VPWR VGND sg13g2_decap_8
XFILLER_5_186 VPWR VGND sg13g2_decap_8
XFILLER_2_893 VPWR VGND sg13g2_decap_8
XFILLER_1_392 VPWR VGND sg13g2_decap_8
XFILLER_37_503 VPWR VGND sg13g2_decap_8
XFILLER_49_385 VPWR VGND sg13g2_decap_8
XFILLER_24_208 VPWR VGND sg13g2_decap_8
XFILLER_21_948 VPWR VGND sg13g2_decap_8
XFILLER_33_775 VPWR VGND sg13g2_decap_8
XFILLER_20_425 VPWR VGND sg13g2_decap_8
XFILLER_32_285 VPWR VGND sg13g2_fill_2
XFILLER_0_819 VPWR VGND sg13g2_decap_8
XFILLER_28_547 VPWR VGND sg13g2_decap_8
XFILLER_15_219 VPWR VGND sg13g2_decap_8
XFILLER_23_230 VPWR VGND sg13g2_decap_8
XFILLER_24_753 VPWR VGND sg13g2_decap_8
XFILLER_11_403 VPWR VGND sg13g2_decap_8
XFILLER_23_11 VPWR VGND sg13g2_decap_8
XFILLER_23_88 VPWR VGND sg13g2_decap_8
XFILLER_20_992 VPWR VGND sg13g2_decap_8
X_060_ VPWR _035_ net47 VGND sg13g2_inv_1
XFILLER_3_613 VPWR VGND sg13g2_decap_8
XFILLER_2_123 VPWR VGND sg13g2_decap_8
XFILLER_47_812 VPWR VGND sg13g2_decap_8
XFILLER_48_63 VPWR VGND sg13g2_decap_8
XFILLER_19_503 VPWR VGND sg13g2_decap_8
XFILLER_46_322 VPWR VGND sg13g2_decap_8
XFILLER_47_889 VPWR VGND sg13g2_decap_8
XFILLER_34_517 VPWR VGND sg13g2_decap_8
XFILLER_46_399 VPWR VGND sg13g2_decap_8
XFILLER_15_742 VPWR VGND sg13g2_decap_8
XFILLER_42_572 VPWR VGND sg13g2_decap_8
XFILLER_30_723 VPWR VGND sg13g2_decap_8
XFILLER_9_46 VPWR VGND sg13g2_decap_8
XFILLER_11_970 VPWR VGND sg13g2_decap_8
XFILLER_10_480 VPWR VGND sg13g2_decap_8
XFILLER_7_952 VPWR VGND sg13g2_decap_8
XFILLER_6_473 VPWR VGND sg13g2_decap_8
XFILLER_9_1026 VPWR VGND sg13g2_fill_2
XFILLER_2_690 VPWR VGND sg13g2_decap_8
XFILLER_49_182 VPWR VGND sg13g2_decap_8
XFILLER_38_834 VPWR VGND sg13g2_decap_8
XFILLER_37_377 VPWR VGND sg13g2_decap_8
XFILLER_40_509 VPWR VGND sg13g2_decap_8
XFILLER_33_572 VPWR VGND sg13g2_decap_8
XFILLER_20_200 VPWR VGND sg13g2_decap_8
XFILLER_21_745 VPWR VGND sg13g2_decap_8
XFILLER_20_277 VPWR VGND sg13g2_decap_8
XFILLER_0_616 VPWR VGND sg13g2_decap_8
XFILLER_48_609 VPWR VGND sg13g2_decap_8
XFILLER_47_119 VPWR VGND sg13g2_decap_8
XFILLER_29_823 VPWR VGND sg13g2_decap_8
XFILLER_18_11 VPWR VGND sg13g2_decap_8
XFILLER_28_300 VPWR VGND sg13g2_decap_8
XFILLER_16_517 VPWR VGND sg13g2_decap_8
XFILLER_18_88 VPWR VGND sg13g2_decap_8
XFILLER_44_859 VPWR VGND sg13g2_decap_8
XFILLER_43_369 VPWR VGND sg13g2_decap_8
XFILLER_24_550 VPWR VGND sg13g2_decap_8
XFILLER_34_54 VPWR VGND sg13g2_decap_8
XFILLER_11_200 VPWR VGND sg13g2_decap_8
XFILLER_12_767 VPWR VGND sg13g2_decap_8
XFILLER_11_277 VPWR VGND sg13g2_decap_8
X_112_ net1 net17 _026_ _027_ VPWR VGND sg13g2_a21o_1
XFILLER_7_259 VPWR VGND sg13g2_decap_8
XFILLER_4_900 VPWR VGND sg13g2_decap_8
XFILLER_3_410 VPWR VGND sg13g2_decap_8
XFILLER_4_977 VPWR VGND sg13g2_decap_8
XFILLER_3_487 VPWR VGND sg13g2_decap_8
XFILLER_1_0 VPWR VGND sg13g2_decap_8
XFILLER_19_311 VPWR VGND sg13g2_decap_8
XFILLER_35_815 VPWR VGND sg13g2_decap_8
XFILLER_47_686 VPWR VGND sg13g2_decap_8
XFILLER_46_196 VPWR VGND sg13g2_decap_8
XFILLER_30_520 VPWR VGND sg13g2_decap_8
XFILLER_30_597 VPWR VGND sg13g2_decap_8
XFILLER_6_270 VPWR VGND sg13g2_decap_8
XFILLER_29_119 VPWR VGND sg13g2_decap_8
XFILLER_38_631 VPWR VGND sg13g2_decap_8
XFILLER_1_91 VPWR VGND sg13g2_decap_8
XFILLER_25_325 VPWR VGND sg13g2_decap_8
XFILLER_26_826 VPWR VGND sg13g2_decap_8
XFILLER_38_1009 VPWR VGND sg13g2_decap_8
XFILLER_34_881 VPWR VGND sg13g2_decap_8
XFILLER_40_306 VPWR VGND sg13g2_decap_8
XFILLER_21_542 VPWR VGND sg13g2_decap_8
XFILLER_4_207 VPWR VGND sg13g2_decap_8
XFILLER_1_903 VPWR VGND sg13g2_decap_8
XFILLER_20_67 VPWR VGND sg13g2_decap_8
XFILLER_0_413 VPWR VGND sg13g2_decap_8
XFILLER_48_406 VPWR VGND sg13g2_decap_8
XFILLER_29_21 VPWR VGND sg13g2_decap_8
XFILLER_29_620 VPWR VGND sg13g2_decap_8
XFILLER_29_98 VPWR VGND sg13g2_decap_8
XFILLER_28_130 VPWR VGND sg13g2_decap_8
XFILLER_17_826 VPWR VGND sg13g2_decap_8
XFILLER_29_697 VPWR VGND sg13g2_decap_8
XFILLER_44_656 VPWR VGND sg13g2_decap_8
XFILLER_45_75 VPWR VGND sg13g2_decap_8
XFILLER_43_166 VPWR VGND sg13g2_decap_8
XFILLER_12_564 VPWR VGND sg13g2_decap_8
XFILLER_40_873 VPWR VGND sg13g2_decap_8
XFILLER_8_557 VPWR VGND sg13g2_decap_8
XFILLER_6_25 VPWR VGND sg13g2_decap_8
XFILLER_4_774 VPWR VGND sg13g2_decap_8
XFILLER_3_284 VPWR VGND sg13g2_decap_8
XFILLER_39_417 VPWR VGND sg13g2_decap_8
XFILLER_0_980 VPWR VGND sg13g2_decap_8
XFILLER_48_973 VPWR VGND sg13g2_decap_8
XFILLER_19_130 VPWR VGND sg13g2_decap_8
XFILLER_47_483 VPWR VGND sg13g2_decap_8
XFILLER_35_612 VPWR VGND sg13g2_decap_8
XFILLER_22_306 VPWR VGND sg13g2_decap_8
XFILLER_34_166 VPWR VGND sg13g2_decap_8
XFILLER_35_689 VPWR VGND sg13g2_decap_8
XFILLER_16_881 VPWR VGND sg13g2_decap_8
XFILLER_31_862 VPWR VGND sg13g2_decap_8
XFILLER_30_394 VPWR VGND sg13g2_decap_8
XFILLER_44_1013 VPWR VGND sg13g2_decap_8
Xheichips25_template_34 VPWR VGND uio_oe[1] sg13g2_tiehi
XFILLER_26_623 VPWR VGND sg13g2_decap_8
XFILLER_39_984 VPWR VGND sg13g2_decap_8
XFILLER_14_829 VPWR VGND sg13g2_decap_8
XFILLER_25_144 VPWR VGND sg13g2_decap_8
XFILLER_15_67 VPWR VGND sg13g2_decap_8
XFILLER_40_158 VPWR VGND sg13g2_decap_8
XFILLER_22_884 VPWR VGND sg13g2_decap_8
XFILLER_31_33 VPWR VGND sg13g2_decap_8
Xoutput22 net27 uo_out[2] VPWR VGND sg13g2_buf_1
XFILLER_1_700 VPWR VGND sg13g2_decap_8
XFILLER_0_210 VPWR VGND sg13g2_decap_8
XFILLER_1_777 VPWR VGND sg13g2_decap_8
XFILLER_48_203 VPWR VGND sg13g2_decap_8
XFILLER_0_287 VPWR VGND sg13g2_decap_8
XFILLER_45_943 VPWR VGND sg13g2_decap_8
XFILLER_17_623 VPWR VGND sg13g2_decap_8
XFILLER_29_494 VPWR VGND sg13g2_decap_8
XFILLER_44_453 VPWR VGND sg13g2_decap_8
XFILLER_16_144 VPWR VGND sg13g2_decap_8
XFILLER_31_103 VPWR VGND sg13g2_decap_8
XFILLER_13_851 VPWR VGND sg13g2_decap_8
XFILLER_9_844 VPWR VGND sg13g2_decap_8
XFILLER_12_361 VPWR VGND sg13g2_decap_8
XFILLER_40_670 VPWR VGND sg13g2_decap_8
XFILLER_8_354 VPWR VGND sg13g2_decap_8
XFILLER_4_571 VPWR VGND sg13g2_decap_8
XFILLER_39_214 VPWR VGND sg13g2_decap_8
XFILLER_48_770 VPWR VGND sg13g2_decap_8
XFILLER_36_921 VPWR VGND sg13g2_decap_8
XFILLER_47_280 VPWR VGND sg13g2_decap_8
XFILLER_36_998 VPWR VGND sg13g2_decap_8
XFILLER_23_648 VPWR VGND sg13g2_decap_8
XFILLER_35_486 VPWR VGND sg13g2_decap_8
XFILLER_30_180 VPWR VGND sg13g2_decap_8
XFILLER_11_1012 VPWR VGND sg13g2_decap_8
XFILLER_2_508 VPWR VGND sg13g2_decap_8
XFILLER_46_707 VPWR VGND sg13g2_decap_8
XFILLER_27_910 VPWR VGND sg13g2_decap_8
XFILLER_39_781 VPWR VGND sg13g2_decap_8
XFILLER_26_11 VPWR VGND sg13g2_decap_8
XFILLER_26_420 VPWR VGND sg13g2_decap_8
XFILLER_38_291 VPWR VGND sg13g2_decap_8
XFILLER_27_987 VPWR VGND sg13g2_decap_8
XFILLER_42_957 VPWR VGND sg13g2_decap_8
XFILLER_14_626 VPWR VGND sg13g2_decap_8
XFILLER_26_88 VPWR VGND sg13g2_decap_8
XFILLER_26_497 VPWR VGND sg13g2_decap_8
XFILLER_41_467 VPWR VGND sg13g2_decap_8
XFILLER_13_158 VPWR VGND sg13g2_decap_8
XFILLER_42_54 VPWR VGND sg13g2_decap_8
XFILLER_22_681 VPWR VGND sg13g2_decap_8
XFILLER_10_865 VPWR VGND sg13g2_decap_8
XFILLER_6_858 VPWR VGND sg13g2_decap_8
XFILLER_5_368 VPWR VGND sg13g2_decap_8
XFILLER_1_574 VPWR VGND sg13g2_decap_8
XFILLER_49_567 VPWR VGND sg13g2_decap_8
XFILLER_18_921 VPWR VGND sg13g2_decap_8
XFILLER_45_740 VPWR VGND sg13g2_decap_8
XFILLER_17_420 VPWR VGND sg13g2_decap_8
XFILLER_44_250 VPWR VGND sg13g2_decap_8
XFILLER_17_497 VPWR VGND sg13g2_decap_8
XFILLER_18_998 VPWR VGND sg13g2_decap_8
XFILLER_20_607 VPWR VGND sg13g2_decap_8
XFILLER_33_957 VPWR VGND sg13g2_decap_8
XFILLER_32_467 VPWR VGND sg13g2_decap_8
XFILLER_9_641 VPWR VGND sg13g2_decap_8
XFILLER_8_151 VPWR VGND sg13g2_decap_8
XFILLER_41_1027 VPWR VGND sg13g2_fill_2
XFILLER_27_217 VPWR VGND sg13g2_decap_8
XFILLER_28_729 VPWR VGND sg13g2_decap_8
XFILLER_24_935 VPWR VGND sg13g2_decap_8
XFILLER_36_795 VPWR VGND sg13g2_decap_8
XFILLER_23_445 VPWR VGND sg13g2_decap_8
XFILLER_12_46 VPWR VGND sg13g2_decap_8
XFILLER_2_305 VPWR VGND sg13g2_decap_8
XFILLER_46_504 VPWR VGND sg13g2_decap_8
XFILLER_37_21 VPWR VGND sg13g2_decap_8
XFILLER_18_228 VPWR VGND sg13g2_fill_1
XFILLER_37_98 VPWR VGND sg13g2_decap_8
XFILLER_14_423 VPWR VGND sg13g2_decap_8
XFILLER_15_924 VPWR VGND sg13g2_decap_8
XFILLER_27_784 VPWR VGND sg13g2_decap_8
XFILLER_42_754 VPWR VGND sg13g2_decap_8
XFILLER_30_905 VPWR VGND sg13g2_decap_8
XFILLER_41_242 VPWR VGND sg13g2_decap_8
XFILLER_10_662 VPWR VGND sg13g2_decap_8
XFILLER_6_655 VPWR VGND sg13g2_decap_8
XFILLER_5_165 VPWR VGND sg13g2_decap_8
XFILLER_2_872 VPWR VGND sg13g2_decap_8
XFILLER_1_371 VPWR VGND sg13g2_decap_8
XFILLER_49_364 VPWR VGND sg13g2_decap_8
XFILLER_37_559 VPWR VGND sg13g2_decap_8
XFILLER_18_795 VPWR VGND sg13g2_decap_8
XFILLER_17_294 VPWR VGND sg13g2_decap_8
XFILLER_33_754 VPWR VGND sg13g2_decap_8
XFILLER_20_404 VPWR VGND sg13g2_decap_8
XFILLER_21_927 VPWR VGND sg13g2_decap_8
XFILLER_32_264 VPWR VGND sg13g2_decap_8
XFILLER_14_990 VPWR VGND sg13g2_decap_8
XFILLER_28_526 VPWR VGND sg13g2_decap_8
XFILLER_24_732 VPWR VGND sg13g2_decap_8
XFILLER_36_592 VPWR VGND sg13g2_decap_8
XFILLER_12_949 VPWR VGND sg13g2_decap_8
XFILLER_11_459 VPWR VGND sg13g2_decap_8
XFILLER_20_971 VPWR VGND sg13g2_decap_8
XFILLER_23_67 VPWR VGND sg13g2_decap_8
XFILLER_2_102 VPWR VGND sg13g2_decap_8
XFILLER_3_669 VPWR VGND sg13g2_decap_8
XFILLER_3_4 VPWR VGND sg13g2_decap_8
XFILLER_2_179 VPWR VGND sg13g2_decap_8
XFILLER_48_42 VPWR VGND sg13g2_decap_8
XFILLER_46_301 VPWR VGND sg13g2_decap_8
XFILLER_47_868 VPWR VGND sg13g2_decap_8
XFILLER_0_49 VPWR VGND sg13g2_decap_8
XFILLER_19_559 VPWR VGND sg13g2_decap_8
XFILLER_46_378 VPWR VGND sg13g2_decap_8
XFILLER_15_721 VPWR VGND sg13g2_decap_8
XFILLER_27_581 VPWR VGND sg13g2_decap_8
XFILLER_42_551 VPWR VGND sg13g2_decap_8
XFILLER_9_25 VPWR VGND sg13g2_decap_8
XFILLER_30_702 VPWR VGND sg13g2_decap_8
XFILLER_14_297 VPWR VGND sg13g2_decap_8
XFILLER_15_798 VPWR VGND sg13g2_decap_8
XFILLER_30_779 VPWR VGND sg13g2_decap_8
XFILLER_7_931 VPWR VGND sg13g2_decap_8
XFILLER_6_452 VPWR VGND sg13g2_decap_8
XFILLER_43_5 VPWR VGND sg13g2_decap_8
XFILLER_9_1005 VPWR VGND sg13g2_decap_8
XFILLER_38_813 VPWR VGND sg13g2_decap_8
XFILLER_49_161 VPWR VGND sg13g2_decap_8
XFILLER_37_356 VPWR VGND sg13g2_decap_8
XFILLER_18_592 VPWR VGND sg13g2_decap_8
XFILLER_33_551 VPWR VGND sg13g2_decap_8
XFILLER_21_724 VPWR VGND sg13g2_decap_8
XFILLER_20_256 VPWR VGND sg13g2_decap_8
XFILLER_47_1022 VPWR VGND sg13g2_decap_8
XFILLER_29_802 VPWR VGND sg13g2_decap_8
XFILLER_18_67 VPWR VGND sg13g2_decap_8
XFILLER_29_879 VPWR VGND sg13g2_decap_8
XFILLER_44_838 VPWR VGND sg13g2_decap_8
XFILLER_28_389 VPWR VGND sg13g2_decap_8
XFILLER_43_348 VPWR VGND sg13g2_decap_8
XFILLER_34_33 VPWR VGND sg13g2_decap_8
XFILLER_12_746 VPWR VGND sg13g2_decap_8
XFILLER_11_256 VPWR VGND sg13g2_decap_8
X_111_ VGND VPWR _026_ net18 net19 sg13g2_or2_1
XFILLER_8_739 VPWR VGND sg13g2_decap_8
XFILLER_7_238 VPWR VGND sg13g2_decap_8
XFILLER_4_956 VPWR VGND sg13g2_decap_8
XFILLER_3_466 VPWR VGND sg13g2_decap_8
XFILLER_38_109 VPWR VGND sg13g2_decap_8
XFILLER_47_665 VPWR VGND sg13g2_decap_8
XFILLER_46_175 VPWR VGND sg13g2_decap_8
XFILLER_19_367 VPWR VGND sg13g2_decap_8
XFILLER_28_890 VPWR VGND sg13g2_decap_8
XFILLER_15_595 VPWR VGND sg13g2_decap_8
XFILLER_30_576 VPWR VGND sg13g2_decap_8
XFILLER_27_0 VPWR VGND sg13g2_decap_8
XFILLER_38_610 VPWR VGND sg13g2_decap_8
XFILLER_26_805 VPWR VGND sg13g2_decap_8
XFILLER_1_70 VPWR VGND sg13g2_decap_8
XFILLER_25_304 VPWR VGND sg13g2_decap_8
XFILLER_38_687 VPWR VGND sg13g2_decap_8
XFILLER_34_860 VPWR VGND sg13g2_decap_8
XFILLER_21_521 VPWR VGND sg13g2_decap_8
XFILLER_33_392 VPWR VGND sg13g2_decap_8
XFILLER_21_598 VPWR VGND sg13g2_decap_8
XFILLER_20_46 VPWR VGND sg13g2_decap_8
XFILLER_1_959 VPWR VGND sg13g2_decap_8
XFILLER_0_469 VPWR VGND sg13g2_decap_8
XFILLER_29_77 VPWR VGND sg13g2_decap_8
XFILLER_17_805 VPWR VGND sg13g2_decap_8
XFILLER_21_1025 VPWR VGND sg13g2_decap_4
XFILLER_29_676 VPWR VGND sg13g2_decap_8
XFILLER_45_54 VPWR VGND sg13g2_decap_8
XFILLER_44_635 VPWR VGND sg13g2_decap_8
XFILLER_16_326 VPWR VGND sg13g2_decap_8
XFILLER_28_197 VPWR VGND sg13g2_decap_8
XFILLER_43_145 VPWR VGND sg13g2_decap_8
XFILLER_12_543 VPWR VGND sg13g2_decap_8
XFILLER_40_852 VPWR VGND sg13g2_decap_8
XFILLER_8_536 VPWR VGND sg13g2_decap_8
XFILLER_4_753 VPWR VGND sg13g2_decap_8
XFILLER_3_263 VPWR VGND sg13g2_decap_8
XFILLER_6_1019 VPWR VGND sg13g2_decap_8
XFILLER_48_952 VPWR VGND sg13g2_decap_8
XFILLER_47_462 VPWR VGND sg13g2_decap_8
XFILLER_19_153 VPWR VGND sg13g2_fill_1
XFILLER_16_860 VPWR VGND sg13g2_decap_8
XFILLER_34_145 VPWR VGND sg13g2_decap_8
XFILLER_35_668 VPWR VGND sg13g2_decap_8
XFILLER_37_1021 VPWR VGND sg13g2_decap_8
XFILLER_15_392 VPWR VGND sg13g2_decap_8
XFILLER_31_841 VPWR VGND sg13g2_decap_8
XFILLER_30_373 VPWR VGND sg13g2_decap_8
Xheichips25_template_35 VPWR VGND uio_oe[2] sg13g2_tiehi
XFILLER_39_963 VPWR VGND sg13g2_decap_8
XFILLER_26_602 VPWR VGND sg13g2_decap_8
XFILLER_25_123 VPWR VGND sg13g2_decap_8
XFILLER_38_484 VPWR VGND sg13g2_decap_8
XFILLER_14_808 VPWR VGND sg13g2_decap_8
XFILLER_26_679 VPWR VGND sg13g2_decap_8
XFILLER_41_649 VPWR VGND sg13g2_decap_8
XFILLER_15_46 VPWR VGND sg13g2_decap_8
XFILLER_25_189 VPWR VGND sg13g2_decap_8
XFILLER_22_863 VPWR VGND sg13g2_decap_8
XFILLER_40_137 VPWR VGND sg13g2_decap_8
XFILLER_21_395 VPWR VGND sg13g2_decap_8
XFILLER_31_12 VPWR VGND sg13g2_decap_8
XFILLER_31_89 VPWR VGND sg13g2_decap_8
Xoutput23 net28 uo_out[3] VPWR VGND sg13g2_buf_1
XFILLER_1_756 VPWR VGND sg13g2_decap_8
XFILLER_49_749 VPWR VGND sg13g2_decap_8
XFILLER_0_266 VPWR VGND sg13g2_decap_8
XFILLER_48_259 VPWR VGND sg13g2_decap_8
XFILLER_45_922 VPWR VGND sg13g2_decap_8
XFILLER_17_602 VPWR VGND sg13g2_decap_8
XFILLER_29_473 VPWR VGND sg13g2_decap_8
XFILLER_44_432 VPWR VGND sg13g2_decap_8
XFILLER_16_123 VPWR VGND sg13g2_decap_8
XFILLER_45_999 VPWR VGND sg13g2_decap_8
XFILLER_17_679 VPWR VGND sg13g2_decap_8
XFILLER_32_649 VPWR VGND sg13g2_decap_8
XFILLER_13_830 VPWR VGND sg13g2_decap_8
XFILLER_31_159 VPWR VGND sg13g2_decap_8
XFILLER_9_823 VPWR VGND sg13g2_decap_8
XFILLER_12_340 VPWR VGND sg13g2_decap_8
XFILLER_8_333 VPWR VGND sg13g2_decap_8
XFILLER_4_550 VPWR VGND sg13g2_decap_8
XFILLER_28_1009 VPWR VGND sg13g2_decap_8
XFILLER_36_900 VPWR VGND sg13g2_decap_8
XFILLER_35_465 VPWR VGND sg13g2_decap_8
XFILLER_36_977 VPWR VGND sg13g2_decap_8
XFILLER_23_627 VPWR VGND sg13g2_decap_8
XFILLER_22_137 VPWR VGND sg13g2_decap_8
XFILLER_7_91 VPWR VGND sg13g2_decap_8
XFILLER_39_760 VPWR VGND sg13g2_decap_8
XFILLER_45_229 VPWR VGND sg13g2_decap_8
XFILLER_38_270 VPWR VGND sg13g2_decap_8
XFILLER_14_605 VPWR VGND sg13g2_decap_8
XFILLER_27_966 VPWR VGND sg13g2_decap_8
XFILLER_42_936 VPWR VGND sg13g2_decap_8
XFILLER_26_67 VPWR VGND sg13g2_decap_8
XFILLER_26_476 VPWR VGND sg13g2_decap_8
XFILLER_41_446 VPWR VGND sg13g2_decap_8
XFILLER_13_137 VPWR VGND sg13g2_decap_8
XFILLER_42_33 VPWR VGND sg13g2_decap_8
XFILLER_22_660 VPWR VGND sg13g2_decap_8
XFILLER_10_844 VPWR VGND sg13g2_decap_8
XFILLER_6_837 VPWR VGND sg13g2_decap_8
XFILLER_5_347 VPWR VGND sg13g2_decap_8
XFILLER_1_553 VPWR VGND sg13g2_decap_8
XFILLER_49_546 VPWR VGND sg13g2_decap_8
XFILLER_18_900 VPWR VGND sg13g2_decap_8
XFILLER_18_977 VPWR VGND sg13g2_decap_8
XFILLER_45_796 VPWR VGND sg13g2_decap_8
XFILLER_17_476 VPWR VGND sg13g2_decap_8
XFILLER_33_936 VPWR VGND sg13g2_decap_8
XFILLER_32_446 VPWR VGND sg13g2_decap_8
XFILLER_9_620 VPWR VGND sg13g2_decap_8
XFILLER_8_130 VPWR VGND sg13g2_decap_8
XFILLER_9_697 VPWR VGND sg13g2_decap_8
XFILLER_41_1006 VPWR VGND sg13g2_decap_8
XFILLER_28_708 VPWR VGND sg13g2_decap_8
XFILLER_24_914 VPWR VGND sg13g2_decap_8
XFILLER_35_262 VPWR VGND sg13g2_decap_4
XFILLER_36_774 VPWR VGND sg13g2_decap_8
XFILLER_23_424 VPWR VGND sg13g2_decap_8
XFILLER_12_25 VPWR VGND sg13g2_decap_8
XFILLER_18_207 VPWR VGND sg13g2_decap_8
XFILLER_15_903 VPWR VGND sg13g2_decap_8
XFILLER_27_763 VPWR VGND sg13g2_decap_8
XFILLER_37_77 VPWR VGND sg13g2_decap_8
XFILLER_14_402 VPWR VGND sg13g2_decap_8
XFILLER_42_733 VPWR VGND sg13g2_decap_8
XFILLER_18_1019 VPWR VGND sg13g2_decap_8
XFILLER_26_295 VPWR VGND sg13g2_fill_2
XFILLER_41_221 VPWR VGND sg13g2_decap_8
XFILLER_14_479 VPWR VGND sg13g2_decap_8
XFILLER_23_991 VPWR VGND sg13g2_decap_8
XFILLER_10_641 VPWR VGND sg13g2_decap_8
XFILLER_6_634 VPWR VGND sg13g2_decap_8
XFILLER_5_144 VPWR VGND sg13g2_decap_8
XFILLER_2_851 VPWR VGND sg13g2_decap_8
XFILLER_1_350 VPWR VGND sg13g2_decap_8
XFILLER_49_343 VPWR VGND sg13g2_decap_8
XFILLER_37_538 VPWR VGND sg13g2_decap_8
XFILLER_17_273 VPWR VGND sg13g2_decap_8
XFILLER_18_774 VPWR VGND sg13g2_decap_8
XFILLER_45_593 VPWR VGND sg13g2_decap_8
XFILLER_33_733 VPWR VGND sg13g2_decap_8
XFILLER_21_906 VPWR VGND sg13g2_decap_8
XFILLER_32_243 VPWR VGND sg13g2_decap_8
XFILLER_9_494 VPWR VGND sg13g2_decap_8
XFILLER_4_81 VPWR VGND sg13g2_decap_8
XFILLER_28_505 VPWR VGND sg13g2_decap_8
XFILLER_24_711 VPWR VGND sg13g2_decap_8
XFILLER_36_571 VPWR VGND sg13g2_decap_8
XFILLER_12_928 VPWR VGND sg13g2_decap_8
XFILLER_24_788 VPWR VGND sg13g2_decap_8
XFILLER_11_438 VPWR VGND sg13g2_decap_8
XFILLER_23_46 VPWR VGND sg13g2_decap_8
XFILLER_23_298 VPWR VGND sg13g2_decap_8
XFILLER_20_950 VPWR VGND sg13g2_decap_8
XFILLER_3_648 VPWR VGND sg13g2_decap_8
XFILLER_2_158 VPWR VGND sg13g2_decap_8
XFILLER_48_21 VPWR VGND sg13g2_decap_8
XFILLER_24_1012 VPWR VGND sg13g2_decap_8
XFILLER_47_847 VPWR VGND sg13g2_decap_8
XFILLER_48_98 VPWR VGND sg13g2_decap_8
XFILLER_19_538 VPWR VGND sg13g2_decap_8
XFILLER_46_357 VPWR VGND sg13g2_decap_8
XFILLER_0_28 VPWR VGND sg13g2_decap_8
XFILLER_15_700 VPWR VGND sg13g2_decap_8
XFILLER_27_560 VPWR VGND sg13g2_decap_8
XFILLER_42_530 VPWR VGND sg13g2_decap_8
XFILLER_14_221 VPWR VGND sg13g2_decap_8
XFILLER_15_777 VPWR VGND sg13g2_decap_8
XFILLER_14_276 VPWR VGND sg13g2_decap_8
XFILLER_7_910 VPWR VGND sg13g2_decap_8
XFILLER_30_758 VPWR VGND sg13g2_decap_8
XFILLER_31_1016 VPWR VGND sg13g2_decap_8
XFILLER_31_1027 VPWR VGND sg13g2_fill_2
XFILLER_6_431 VPWR VGND sg13g2_decap_8
XFILLER_7_987 VPWR VGND sg13g2_decap_8
XFILLER_9_1028 VPWR VGND sg13g2_fill_1
XFILLER_36_5 VPWR VGND sg13g2_decap_8
XFILLER_49_140 VPWR VGND sg13g2_decap_8
XFILLER_37_313 VPWR VGND sg13g2_decap_4
XFILLER_37_335 VPWR VGND sg13g2_decap_8
XFILLER_38_869 VPWR VGND sg13g2_decap_8
XFILLER_18_571 VPWR VGND sg13g2_decap_8
XFILLER_45_390 VPWR VGND sg13g2_decap_8
XFILLER_33_530 VPWR VGND sg13g2_decap_8
XFILLER_21_703 VPWR VGND sg13g2_decap_8
XFILLER_20_235 VPWR VGND sg13g2_decap_8
XFILLER_9_291 VPWR VGND sg13g2_decap_8
XFILLER_47_1001 VPWR VGND sg13g2_decap_8
XFILLER_18_46 VPWR VGND sg13g2_decap_8
XFILLER_28_335 VPWR VGND sg13g2_decap_8
XFILLER_28_346 VPWR VGND sg13g2_fill_2
XFILLER_29_858 VPWR VGND sg13g2_decap_8
XFILLER_44_817 VPWR VGND sg13g2_decap_8
XFILLER_28_368 VPWR VGND sg13g2_decap_8
XFILLER_43_327 VPWR VGND sg13g2_decap_8
XFILLER_34_12 VPWR VGND sg13g2_decap_8
XFILLER_12_725 VPWR VGND sg13g2_decap_8
XFILLER_24_585 VPWR VGND sg13g2_decap_8
XFILLER_34_89 VPWR VGND sg13g2_decap_8
XFILLER_8_718 VPWR VGND sg13g2_decap_8
XFILLER_11_235 VPWR VGND sg13g2_decap_8
X_110_ net18 _024_ net19 _025_ VPWR VGND sg13g2_nand3_1
XFILLER_7_217 VPWR VGND sg13g2_decap_8
Xclkload0 clknet_2_0__leaf_clk clkload0/X VPWR VGND sg13g2_buf_1
XFILLER_4_935 VPWR VGND sg13g2_decap_8
XFILLER_3_445 VPWR VGND sg13g2_decap_8
XFILLER_47_644 VPWR VGND sg13g2_decap_8
XFILLER_19_346 VPWR VGND sg13g2_decap_8
XFILLER_46_154 VPWR VGND sg13g2_decap_8
XFILLER_34_338 VPWR VGND sg13g2_decap_8
XFILLER_43_894 VPWR VGND sg13g2_decap_8
XFILLER_15_574 VPWR VGND sg13g2_decap_8
XFILLER_30_555 VPWR VGND sg13g2_decap_8
XFILLER_7_784 VPWR VGND sg13g2_decap_8
XFILLER_38_666 VPWR VGND sg13g2_decap_8
XFILLER_37_187 VPWR VGND sg13g2_decap_8
XFILLER_21_500 VPWR VGND sg13g2_decap_8
XFILLER_33_371 VPWR VGND sg13g2_decap_8
XFILLER_14_1011 VPWR VGND sg13g2_decap_8
XFILLER_21_577 VPWR VGND sg13g2_decap_8
XFILLER_20_25 VPWR VGND sg13g2_decap_8
XFILLER_1_938 VPWR VGND sg13g2_decap_8
XFILLER_0_448 VPWR VGND sg13g2_decap_8
XFILLER_29_56 VPWR VGND sg13g2_decap_8
XFILLER_21_1004 VPWR VGND sg13g2_decap_8
XFILLER_29_655 VPWR VGND sg13g2_decap_8
XFILLER_44_614 VPWR VGND sg13g2_decap_8
XFILLER_16_305 VPWR VGND sg13g2_decap_8
XFILLER_45_33 VPWR VGND sg13g2_decap_8
XFILLER_43_124 VPWR VGND sg13g2_decap_8
XFILLER_16_349 VPWR VGND sg13g2_decap_8
XFILLER_28_176 VPWR VGND sg13g2_decap_8
XFILLER_25_894 VPWR VGND sg13g2_decap_8
XFILLER_12_522 VPWR VGND sg13g2_decap_8
XFILLER_24_393 VPWR VGND sg13g2_decap_4
XFILLER_40_831 VPWR VGND sg13g2_decap_8
XFILLER_8_515 VPWR VGND sg13g2_decap_8
XFILLER_12_599 VPWR VGND sg13g2_decap_8
XFILLER_4_732 VPWR VGND sg13g2_decap_8
XFILLER_3_242 VPWR VGND sg13g2_decap_8
XFILLER_48_931 VPWR VGND sg13g2_decap_8
XFILLER_47_441 VPWR VGND sg13g2_decap_8
XFILLER_34_124 VPWR VGND sg13g2_decap_8
XFILLER_35_647 VPWR VGND sg13g2_decap_8
XFILLER_23_809 VPWR VGND sg13g2_decap_8
XFILLER_37_1000 VPWR VGND sg13g2_decap_8
XFILLER_15_371 VPWR VGND sg13g2_decap_8
XFILLER_31_820 VPWR VGND sg13g2_decap_8
XFILLER_43_691 VPWR VGND sg13g2_decap_8
XFILLER_30_352 VPWR VGND sg13g2_decap_8
XFILLER_31_897 VPWR VGND sg13g2_decap_8
XFILLER_7_581 VPWR VGND sg13g2_decap_8
Xheichips25_template_36 VPWR VGND uio_oe[3] sg13g2_tiehi
XFILLER_39_942 VPWR VGND sg13g2_decap_8
XFILLER_38_463 VPWR VGND sg13g2_decap_8
XFILLER_25_102 VPWR VGND sg13g2_decap_8
XFILLER_26_658 VPWR VGND sg13g2_decap_8
XFILLER_41_628 VPWR VGND sg13g2_decap_8
XFILLER_13_319 VPWR VGND sg13g2_decap_8
XFILLER_15_25 VPWR VGND sg13g2_decap_8
XFILLER_25_168 VPWR VGND sg13g2_decap_8
XFILLER_40_116 VPWR VGND sg13g2_decap_8
XFILLER_22_842 VPWR VGND sg13g2_decap_8
XFILLER_21_374 VPWR VGND sg13g2_decap_8
XFILLER_5_529 VPWR VGND sg13g2_decap_8
XFILLER_31_68 VPWR VGND sg13g2_decap_8
Xoutput24 net29 uo_out[4] VPWR VGND sg13g2_buf_1
XFILLER_1_735 VPWR VGND sg13g2_decap_8
XFILLER_0_245 VPWR VGND sg13g2_decap_8
XFILLER_49_728 VPWR VGND sg13g2_decap_8
XFILLER_48_238 VPWR VGND sg13g2_decap_8
XFILLER_45_901 VPWR VGND sg13g2_decap_8
XFILLER_29_452 VPWR VGND sg13g2_decap_8
XFILLER_44_411 VPWR VGND sg13g2_decap_8
XFILLER_16_102 VPWR VGND sg13g2_decap_8
XFILLER_45_978 VPWR VGND sg13g2_decap_8
XFILLER_17_658 VPWR VGND sg13g2_decap_8
XFILLER_44_488 VPWR VGND sg13g2_decap_8
XFILLER_16_179 VPWR VGND sg13g2_decap_8
XFILLER_32_628 VPWR VGND sg13g2_decap_8
XFILLER_9_802 VPWR VGND sg13g2_decap_8
XFILLER_25_691 VPWR VGND sg13g2_decap_8
XFILLER_31_138 VPWR VGND sg13g2_decap_8
XFILLER_8_312 VPWR VGND sg13g2_decap_8
XFILLER_13_886 VPWR VGND sg13g2_decap_8
XFILLER_12_396 VPWR VGND sg13g2_decap_8
XFILLER_9_879 VPWR VGND sg13g2_decap_8
XFILLER_8_389 VPWR VGND sg13g2_decap_8
XFILLER_39_249 VPWR VGND sg13g2_decap_8
XFILLER_11_4 VPWR VGND sg13g2_decap_8
XFILLER_36_956 VPWR VGND sg13g2_decap_8
XFILLER_23_606 VPWR VGND sg13g2_decap_8
XFILLER_35_444 VPWR VGND sg13g2_decap_8
XFILLER_22_116 VPWR VGND sg13g2_decap_8
XFILLER_31_694 VPWR VGND sg13g2_decap_8
XFILLER_7_70 VPWR VGND sg13g2_decap_8
XFILLER_45_208 VPWR VGND sg13g2_decap_8
XFILLER_27_945 VPWR VGND sg13g2_decap_8
XFILLER_26_46 VPWR VGND sg13g2_decap_8
XFILLER_26_455 VPWR VGND sg13g2_decap_8
XFILLER_42_915 VPWR VGND sg13g2_decap_8
XFILLER_41_425 VPWR VGND sg13g2_decap_8
XFILLER_13_116 VPWR VGND sg13g2_decap_8
XFILLER_42_12 VPWR VGND sg13g2_decap_8
XFILLER_9_109 VPWR VGND sg13g2_decap_8
XFILLER_10_823 VPWR VGND sg13g2_decap_8
XFILLER_42_89 VPWR VGND sg13g2_decap_8
XFILLER_6_816 VPWR VGND sg13g2_decap_8
XFILLER_5_326 VPWR VGND sg13g2_decap_8
XFILLER_1_532 VPWR VGND sg13g2_decap_8
XFILLER_3_39 VPWR VGND sg13g2_decap_8
XFILLER_49_525 VPWR VGND sg13g2_decap_8
XFILLER_36_208 VPWR VGND sg13g2_decap_8
XFILLER_29_271 VPWR VGND sg13g2_decap_8
XFILLER_17_455 VPWR VGND sg13g2_decap_8
XFILLER_18_956 VPWR VGND sg13g2_decap_8
XFILLER_45_775 VPWR VGND sg13g2_decap_8
XFILLER_33_915 VPWR VGND sg13g2_decap_8
XFILLER_44_285 VPWR VGND sg13g2_decap_8
XFILLER_32_425 VPWR VGND sg13g2_decap_8
XFILLER_34_1014 VPWR VGND sg13g2_decap_8
XFILLER_41_992 VPWR VGND sg13g2_decap_8
XFILLER_13_683 VPWR VGND sg13g2_decap_8
XFILLER_9_676 VPWR VGND sg13g2_decap_8
XFILLER_12_193 VPWR VGND sg13g2_decap_8
XFILLER_8_186 VPWR VGND sg13g2_decap_8
XFILLER_5_893 VPWR VGND sg13g2_decap_8
XFILLER_36_753 VPWR VGND sg13g2_decap_8
XFILLER_23_403 VPWR VGND sg13g2_decap_8
XFILLER_35_241 VPWR VGND sg13g2_decap_8
XFILLER_35_285 VPWR VGND sg13g2_decap_8
XFILLER_35_296 VPWR VGND sg13g2_fill_2
XFILLER_32_992 VPWR VGND sg13g2_decap_8
XFILLER_31_491 VPWR VGND sg13g2_decap_8
XFILLER_46_539 VPWR VGND sg13g2_decap_8
XFILLER_2_1012 VPWR VGND sg13g2_decap_8
XFILLER_37_56 VPWR VGND sg13g2_decap_8
XFILLER_27_742 VPWR VGND sg13g2_decap_8
XFILLER_42_712 VPWR VGND sg13g2_decap_8
XFILLER_15_959 VPWR VGND sg13g2_decap_8
XFILLER_26_274 VPWR VGND sg13g2_decap_8
XFILLER_41_200 VPWR VGND sg13g2_decap_8
XFILLER_42_789 VPWR VGND sg13g2_decap_8
XFILLER_14_458 VPWR VGND sg13g2_decap_8
XFILLER_23_970 VPWR VGND sg13g2_decap_8
XFILLER_41_299 VPWR VGND sg13g2_decap_8
XFILLER_41_277 VPWR VGND sg13g2_fill_2
XFILLER_10_620 VPWR VGND sg13g2_decap_8
XFILLER_6_613 VPWR VGND sg13g2_decap_8
XFILLER_10_697 VPWR VGND sg13g2_decap_8
XFILLER_5_123 VPWR VGND sg13g2_decap_8
XFILLER_2_830 VPWR VGND sg13g2_decap_8
XFILLER_49_322 VPWR VGND sg13g2_decap_8
XFILLER_49_399 VPWR VGND sg13g2_decap_8
XFILLER_37_517 VPWR VGND sg13g2_decap_8
XFILLER_18_753 VPWR VGND sg13g2_decap_8
XFILLER_45_572 VPWR VGND sg13g2_decap_8
XFILLER_17_252 VPWR VGND sg13g2_decap_8
XFILLER_33_712 VPWR VGND sg13g2_decap_8
XFILLER_32_222 VPWR VGND sg13g2_decap_8
XFILLER_33_789 VPWR VGND sg13g2_decap_8
XFILLER_20_439 VPWR VGND sg13g2_decap_8
XFILLER_32_299 VPWR VGND sg13g2_decap_8
XFILLER_13_480 VPWR VGND sg13g2_decap_8
XFILLER_9_473 VPWR VGND sg13g2_decap_8
XFILLER_5_690 VPWR VGND sg13g2_decap_8
XFILLER_4_60 VPWR VGND sg13g2_decap_8
XFILLER_43_509 VPWR VGND sg13g2_decap_8
XFILLER_36_550 VPWR VGND sg13g2_decap_8
XFILLER_23_211 VPWR VGND sg13g2_decap_8
XFILLER_23_222 VPWR VGND sg13g2_fill_2
XFILLER_12_907 VPWR VGND sg13g2_decap_8
XFILLER_23_244 VPWR VGND sg13g2_decap_8
XFILLER_24_767 VPWR VGND sg13g2_decap_8
XFILLER_11_417 VPWR VGND sg13g2_decap_8
XFILLER_23_25 VPWR VGND sg13g2_decap_8
XFILLER_23_288 VPWR VGND sg13g2_fill_1
XFILLER_3_627 VPWR VGND sg13g2_decap_8
XFILLER_2_137 VPWR VGND sg13g2_decap_8
XFILLER_47_826 VPWR VGND sg13g2_decap_8
XFILLER_48_77 VPWR VGND sg13g2_decap_8
XFILLER_19_517 VPWR VGND sg13g2_decap_8
XFILLER_46_336 VPWR VGND sg13g2_decap_8
XFILLER_14_200 VPWR VGND sg13g2_decap_8
XFILLER_14_255 VPWR VGND sg13g2_decap_8
XFILLER_15_756 VPWR VGND sg13g2_decap_8
XFILLER_42_586 VPWR VGND sg13g2_decap_8
XFILLER_30_737 VPWR VGND sg13g2_decap_8
XFILLER_6_410 VPWR VGND sg13g2_decap_8
XFILLER_11_984 VPWR VGND sg13g2_decap_8
XFILLER_10_494 VPWR VGND sg13g2_decap_8
XFILLER_7_966 VPWR VGND sg13g2_decap_8
XFILLER_6_487 VPWR VGND sg13g2_decap_8
XFILLER_38_848 VPWR VGND sg13g2_decap_8
XFILLER_49_196 VPWR VGND sg13g2_decap_8
XFILLER_18_550 VPWR VGND sg13g2_decap_8
XFILLER_25_509 VPWR VGND sg13g2_decap_8
XFILLER_20_214 VPWR VGND sg13g2_decap_8
XFILLER_33_586 VPWR VGND sg13g2_decap_8
XFILLER_21_759 VPWR VGND sg13g2_decap_8
XFILLER_9_270 VPWR VGND sg13g2_decap_8
XFILLER_18_25 VPWR VGND sg13g2_decap_8
XFILLER_28_314 VPWR VGND sg13g2_decap_8
XFILLER_29_837 VPWR VGND sg13g2_decap_8
XFILLER_43_306 VPWR VGND sg13g2_decap_8
XFILLER_37_881 VPWR VGND sg13g2_decap_8
XFILLER_12_704 VPWR VGND sg13g2_decap_8
XFILLER_24_564 VPWR VGND sg13g2_decap_8
XFILLER_11_214 VPWR VGND sg13g2_decap_8
XFILLER_34_68 VPWR VGND sg13g2_decap_8
Xclkload1 clknet_2_1__leaf_clk clkload1/X VPWR VGND sg13g2_buf_1
XFILLER_4_914 VPWR VGND sg13g2_decap_8
XFILLER_3_424 VPWR VGND sg13g2_decap_8
XFILLER_47_623 VPWR VGND sg13g2_decap_8
XFILLER_46_133 VPWR VGND sg13g2_decap_8
XFILLER_19_325 VPWR VGND sg13g2_decap_8
XFILLER_35_829 VPWR VGND sg13g2_decap_8
XFILLER_34_317 VPWR VGND sg13g2_decap_8
XFILLER_15_553 VPWR VGND sg13g2_decap_8
XFILLER_43_873 VPWR VGND sg13g2_decap_8
XFILLER_42_383 VPWR VGND sg13g2_decap_8
XFILLER_30_534 VPWR VGND sg13g2_decap_8
XFILLER_11_781 VPWR VGND sg13g2_decap_8
XFILLER_10_291 VPWR VGND sg13g2_decap_8
XFILLER_7_763 VPWR VGND sg13g2_decap_8
XFILLER_6_284 VPWR VGND sg13g2_decap_8
XFILLER_41_4 VPWR VGND sg13g2_decap_8
XFILLER_3_991 VPWR VGND sg13g2_decap_8
XFILLER_37_133 VPWR VGND sg13g2_decap_8
XFILLER_38_645 VPWR VGND sg13g2_decap_8
XFILLER_19_881 VPWR VGND sg13g2_decap_8
XFILLER_25_339 VPWR VGND sg13g2_decap_8
XFILLER_34_895 VPWR VGND sg13g2_decap_8
XFILLER_21_556 VPWR VGND sg13g2_decap_8
XFILLER_1_917 VPWR VGND sg13g2_decap_8
XFILLER_0_427 VPWR VGND sg13g2_decap_8
XFILLER_29_35 VPWR VGND sg13g2_decap_8
XFILLER_29_634 VPWR VGND sg13g2_decap_8
XFILLER_45_12 VPWR VGND sg13g2_decap_8
XFILLER_28_144 VPWR VGND sg13g2_decap_4
XFILLER_43_103 VPWR VGND sg13g2_decap_8
XFILLER_45_89 VPWR VGND sg13g2_decap_8
XFILLER_12_501 VPWR VGND sg13g2_decap_8
XFILLER_24_372 VPWR VGND sg13g2_decap_4
XFILLER_25_873 VPWR VGND sg13g2_decap_8
XFILLER_31_309 VPWR VGND sg13g2_decap_8
XFILLER_40_810 VPWR VGND sg13g2_decap_8
XFILLER_12_578 VPWR VGND sg13g2_decap_8
XFILLER_40_887 VPWR VGND sg13g2_decap_8
XFILLER_6_39 VPWR VGND sg13g2_decap_8
XFILLER_4_711 VPWR VGND sg13g2_decap_8
XFILLER_3_221 VPWR VGND sg13g2_decap_8
XFILLER_10_81 VPWR VGND sg13g2_decap_8
XFILLER_4_788 VPWR VGND sg13g2_decap_8
XFILLER_3_298 VPWR VGND sg13g2_decap_8
XFILLER_48_910 VPWR VGND sg13g2_decap_8
XFILLER_47_420 VPWR VGND sg13g2_decap_8
XFILLER_0_994 VPWR VGND sg13g2_decap_8
XFILLER_48_987 VPWR VGND sg13g2_decap_8
XFILLER_19_144 VPWR VGND sg13g2_decap_8
XFILLER_47_497 VPWR VGND sg13g2_decap_8
XFILLER_19_199 VPWR VGND sg13g2_decap_8
XFILLER_34_103 VPWR VGND sg13g2_decap_8
XFILLER_35_626 VPWR VGND sg13g2_decap_8
XFILLER_43_670 VPWR VGND sg13g2_decap_8
XFILLER_15_350 VPWR VGND sg13g2_decap_8
XFILLER_16_895 VPWR VGND sg13g2_decap_8
XFILLER_42_180 VPWR VGND sg13g2_decap_8
XFILLER_31_876 VPWR VGND sg13g2_decap_8
XFILLER_7_560 VPWR VGND sg13g2_decap_8
XFILLER_44_1027 VPWR VGND sg13g2_fill_2
XFILLER_39_921 VPWR VGND sg13g2_decap_8
Xheichips25_template_37 VPWR VGND uio_oe[4] sg13g2_tiehi
XFILLER_38_442 VPWR VGND sg13g2_decap_8
XFILLER_26_637 VPWR VGND sg13g2_decap_8
XFILLER_39_998 VPWR VGND sg13g2_decap_8
XFILLER_41_607 VPWR VGND sg13g2_decap_8
XFILLER_22_821 VPWR VGND sg13g2_decap_8
XFILLER_34_692 VPWR VGND sg13g2_decap_8
XFILLER_21_353 VPWR VGND sg13g2_decap_8
XFILLER_22_898 VPWR VGND sg13g2_decap_8
XFILLER_5_508 VPWR VGND sg13g2_decap_8
XFILLER_31_47 VPWR VGND sg13g2_decap_8
Xoutput25 net30 uo_out[5] VPWR VGND sg13g2_buf_1
XFILLER_1_714 VPWR VGND sg13g2_decap_8
XFILLER_49_707 VPWR VGND sg13g2_decap_8
XFILLER_0_224 VPWR VGND sg13g2_decap_8
XFILLER_48_217 VPWR VGND sg13g2_decap_8
XFILLER_29_431 VPWR VGND sg13g2_decap_8
XFILLER_17_637 VPWR VGND sg13g2_decap_8
XFILLER_45_957 VPWR VGND sg13g2_decap_8
XFILLER_44_467 VPWR VGND sg13g2_decap_8
XFILLER_16_158 VPWR VGND sg13g2_decap_8
XFILLER_25_670 VPWR VGND sg13g2_decap_8
XFILLER_32_607 VPWR VGND sg13g2_decap_8
XFILLER_31_117 VPWR VGND sg13g2_decap_8
XFILLER_13_865 VPWR VGND sg13g2_decap_8
XFILLER_9_858 VPWR VGND sg13g2_decap_8
XFILLER_12_375 VPWR VGND sg13g2_decap_8
XFILLER_40_684 VPWR VGND sg13g2_decap_8
XFILLER_8_368 VPWR VGND sg13g2_decap_8
XFILLER_4_585 VPWR VGND sg13g2_decap_8
XFILLER_0_791 VPWR VGND sg13g2_decap_8
XFILLER_39_228 VPWR VGND sg13g2_decap_8
XFILLER_48_784 VPWR VGND sg13g2_decap_8
XFILLER_35_423 VPWR VGND sg13g2_decap_8
XFILLER_36_935 VPWR VGND sg13g2_decap_8
XFILLER_47_294 VPWR VGND sg13g2_decap_8
XFILLER_16_692 VPWR VGND sg13g2_decap_8
XFILLER_31_673 VPWR VGND sg13g2_decap_8
XFILLER_30_194 VPWR VGND sg13g2_decap_8
XFILLER_11_1026 VPWR VGND sg13g2_fill_2
XFILLER_27_924 VPWR VGND sg13g2_decap_8
XFILLER_39_795 VPWR VGND sg13g2_decap_8
XFILLER_26_25 VPWR VGND sg13g2_decap_8
XFILLER_26_434 VPWR VGND sg13g2_decap_8
XFILLER_41_404 VPWR VGND sg13g2_decap_8
XFILLER_35_990 VPWR VGND sg13g2_decap_8
XFILLER_10_802 VPWR VGND sg13g2_decap_8
XFILLER_42_68 VPWR VGND sg13g2_decap_8
XFILLER_22_695 VPWR VGND sg13g2_decap_8
XFILLER_10_879 VPWR VGND sg13g2_decap_8
XFILLER_21_183 VPWR VGND sg13g2_decap_8
XFILLER_5_305 VPWR VGND sg13g2_decap_8
XFILLER_1_511 VPWR VGND sg13g2_decap_8
XFILLER_3_18 VPWR VGND sg13g2_decap_8
XFILLER_49_504 VPWR VGND sg13g2_decap_8
XFILLER_27_1022 VPWR VGND sg13g2_decap_8
XFILLER_1_588 VPWR VGND sg13g2_decap_8
XFILLER_18_935 VPWR VGND sg13g2_decap_8
XFILLER_29_250 VPWR VGND sg13g2_decap_8
XFILLER_45_754 VPWR VGND sg13g2_decap_8
XFILLER_17_434 VPWR VGND sg13g2_decap_8
XFILLER_44_264 VPWR VGND sg13g2_decap_8
XFILLER_32_404 VPWR VGND sg13g2_decap_8
XFILLER_41_971 VPWR VGND sg13g2_decap_8
XFILLER_13_662 VPWR VGND sg13g2_decap_8
XFILLER_12_172 VPWR VGND sg13g2_decap_8
XFILLER_40_481 VPWR VGND sg13g2_decap_8
XFILLER_9_655 VPWR VGND sg13g2_decap_8
XFILLER_8_165 VPWR VGND sg13g2_decap_8
XFILLER_5_872 VPWR VGND sg13g2_decap_8
XFILLER_4_382 VPWR VGND sg13g2_decap_8
XFILLER_48_581 VPWR VGND sg13g2_decap_8
XFILLER_36_732 VPWR VGND sg13g2_decap_8
XFILLER_24_949 VPWR VGND sg13g2_decap_8
XFILLER_23_459 VPWR VGND sg13g2_decap_8
XFILLER_10_109 VPWR VGND sg13g2_decap_8
XFILLER_31_470 VPWR VGND sg13g2_decap_8
XFILLER_32_971 VPWR VGND sg13g2_decap_8
XFILLER_3_809 VPWR VGND sg13g2_decap_8
XFILLER_2_319 VPWR VGND sg13g2_decap_8
XFILLER_46_518 VPWR VGND sg13g2_decap_8
XFILLER_27_721 VPWR VGND sg13g2_decap_8
XFILLER_37_35 VPWR VGND sg13g2_decap_8
XFILLER_39_592 VPWR VGND sg13g2_decap_8
XFILLER_26_253 VPWR VGND sg13g2_decap_8
XFILLER_14_437 VPWR VGND sg13g2_decap_8
XFILLER_15_938 VPWR VGND sg13g2_decap_8
XFILLER_27_798 VPWR VGND sg13g2_decap_8
XFILLER_42_768 VPWR VGND sg13g2_decap_8
XFILLER_30_919 VPWR VGND sg13g2_decap_8
XFILLER_41_256 VPWR VGND sg13g2_decap_8
XFILLER_22_492 VPWR VGND sg13g2_decap_8
XFILLER_10_676 VPWR VGND sg13g2_decap_8
XFILLER_5_102 VPWR VGND sg13g2_decap_8
XFILLER_6_669 VPWR VGND sg13g2_decap_8
XFILLER_5_179 VPWR VGND sg13g2_decap_8
XFILLER_49_301 VPWR VGND sg13g2_decap_8
XFILLER_2_886 VPWR VGND sg13g2_decap_8
XFILLER_1_385 VPWR VGND sg13g2_decap_8
XFILLER_49_378 VPWR VGND sg13g2_decap_8
XFILLER_18_732 VPWR VGND sg13g2_decap_8
XFILLER_45_551 VPWR VGND sg13g2_decap_8
XFILLER_17_231 VPWR VGND sg13g2_decap_8
XFILLER_32_201 VPWR VGND sg13g2_decap_8
XFILLER_33_768 VPWR VGND sg13g2_decap_8
XFILLER_20_418 VPWR VGND sg13g2_decap_8
XFILLER_32_278 VPWR VGND sg13g2_decap_8
XFILLER_9_452 VPWR VGND sg13g2_decap_8
XFILLER_24_746 VPWR VGND sg13g2_decap_8
XFILLER_20_985 VPWR VGND sg13g2_decap_8
XFILLER_3_606 VPWR VGND sg13g2_decap_8
XFILLER_2_116 VPWR VGND sg13g2_decap_8
XFILLER_47_805 VPWR VGND sg13g2_decap_8
XFILLER_48_56 VPWR VGND sg13g2_decap_8
XFILLER_46_315 VPWR VGND sg13g2_decap_8
XFILLER_15_735 VPWR VGND sg13g2_decap_8
XFILLER_27_595 VPWR VGND sg13g2_decap_8
XFILLER_42_565 VPWR VGND sg13g2_decap_8
XFILLER_9_39 VPWR VGND sg13g2_decap_8
XFILLER_30_716 VPWR VGND sg13g2_decap_8
XFILLER_11_963 VPWR VGND sg13g2_decap_8
XFILLER_10_473 VPWR VGND sg13g2_decap_8
XFILLER_7_945 VPWR VGND sg13g2_decap_8
XFILLER_13_81 VPWR VGND sg13g2_decap_8
XFILLER_6_466 VPWR VGND sg13g2_decap_8
XFILLER_9_1019 VPWR VGND sg13g2_decap_8
XFILLER_2_683 VPWR VGND sg13g2_decap_8
XFILLER_1_182 VPWR VGND sg13g2_decap_8
XFILLER_49_175 VPWR VGND sg13g2_decap_8
XFILLER_38_827 VPWR VGND sg13g2_decap_8
XFILLER_46_882 VPWR VGND sg13g2_decap_8
XFILLER_21_738 VPWR VGND sg13g2_decap_8
XFILLER_33_565 VPWR VGND sg13g2_decap_8
XFILLER_0_609 VPWR VGND sg13g2_decap_8
XFILLER_29_816 VPWR VGND sg13g2_decap_8
XFILLER_37_860 VPWR VGND sg13g2_decap_8
XFILLER_24_543 VPWR VGND sg13g2_decap_8
XFILLER_34_47 VPWR VGND sg13g2_decap_8
Xclkload2 clknet_2_3__leaf_clk clkload2/X VPWR VGND sg13g2_buf_1
XFILLER_20_782 VPWR VGND sg13g2_decap_8
XFILLER_3_403 VPWR VGND sg13g2_decap_8
XFILLER_47_602 VPWR VGND sg13g2_decap_8
XFILLER_19_304 VPWR VGND sg13g2_decap_8
XFILLER_46_112 VPWR VGND sg13g2_decap_8
XFILLER_47_679 VPWR VGND sg13g2_decap_8
XFILLER_35_808 VPWR VGND sg13g2_decap_8
XFILLER_46_189 VPWR VGND sg13g2_decap_8
XFILLER_43_852 VPWR VGND sg13g2_decap_8
XFILLER_15_532 VPWR VGND sg13g2_decap_8
XFILLER_27_392 VPWR VGND sg13g2_decap_8
XFILLER_42_362 VPWR VGND sg13g2_decap_8
XFILLER_30_513 VPWR VGND sg13g2_decap_8
XFILLER_11_760 VPWR VGND sg13g2_decap_8
XFILLER_10_270 VPWR VGND sg13g2_decap_8
XFILLER_7_742 VPWR VGND sg13g2_decap_8
XFILLER_6_263 VPWR VGND sg13g2_decap_8
X_099_ net2 net3 mod1.qam16_mod.q_level\[2\] VPWR VGND sg13g2_xor2_1
XFILLER_3_970 VPWR VGND sg13g2_decap_8
XFILLER_2_480 VPWR VGND sg13g2_decap_8
XFILLER_37_112 VPWR VGND sg13g2_decap_8
XFILLER_38_624 VPWR VGND sg13g2_decap_8
XFILLER_19_860 VPWR VGND sg13g2_decap_8
XFILLER_26_819 VPWR VGND sg13g2_decap_8
XFILLER_1_84 VPWR VGND sg13g2_decap_8
XFILLER_25_318 VPWR VGND sg13g2_decap_8
XFILLER_33_340 VPWR VGND sg13g2_decap_8
XFILLER_34_874 VPWR VGND sg13g2_decap_8
XFILLER_21_535 VPWR VGND sg13g2_decap_8
XFILLER_0_406 VPWR VGND sg13g2_decap_8
XFILLER_29_14 VPWR VGND sg13g2_decap_8
XFILLER_29_613 VPWR VGND sg13g2_decap_8
XFILLER_28_123 VPWR VGND sg13g2_decap_8
XFILLER_17_819 VPWR VGND sg13g2_decap_8
XFILLER_44_649 VPWR VGND sg13g2_decap_8
XFILLER_45_68 VPWR VGND sg13g2_decap_8
XFILLER_43_159 VPWR VGND sg13g2_decap_8
XFILLER_25_852 VPWR VGND sg13g2_decap_8
XFILLER_24_351 VPWR VGND sg13g2_decap_8
XFILLER_12_557 VPWR VGND sg13g2_decap_8
XFILLER_40_866 VPWR VGND sg13g2_decap_8
XFILLER_6_18 VPWR VGND sg13g2_decap_8
XFILLER_3_200 VPWR VGND sg13g2_decap_8
XFILLER_4_767 VPWR VGND sg13g2_decap_8
XFILLER_10_60 VPWR VGND sg13g2_decap_8
XFILLER_3_277 VPWR VGND sg13g2_decap_8
XFILLER_0_973 VPWR VGND sg13g2_decap_8
XFILLER_19_123 VPWR VGND sg13g2_decap_8
XFILLER_48_966 VPWR VGND sg13g2_decap_8
XFILLER_35_605 VPWR VGND sg13g2_decap_8
XFILLER_47_476 VPWR VGND sg13g2_decap_8
XFILLER_16_874 VPWR VGND sg13g2_decap_8
XFILLER_34_159 VPWR VGND sg13g2_decap_8
XFILLER_31_855 VPWR VGND sg13g2_decap_8
XFILLER_30_332 VPWR VGND sg13g2_fill_2
XFILLER_30_387 VPWR VGND sg13g2_decap_8
XFILLER_44_1006 VPWR VGND sg13g2_decap_8
XFILLER_39_900 VPWR VGND sg13g2_decap_8
XFILLER_38_421 VPWR VGND sg13g2_decap_8
Xheichips25_template_38 VPWR VGND uio_oe[5] sg13g2_tiehi
XFILLER_39_977 VPWR VGND sg13g2_decap_8
XFILLER_26_616 VPWR VGND sg13g2_decap_8
XFILLER_38_498 VPWR VGND sg13g2_decap_8
XFILLER_25_137 VPWR VGND sg13g2_decap_8
XFILLER_22_800 VPWR VGND sg13g2_decap_8
XFILLER_34_671 VPWR VGND sg13g2_decap_8
XFILLER_22_877 VPWR VGND sg13g2_decap_8
XFILLER_31_26 VPWR VGND sg13g2_decap_8
Xoutput26 net31 uo_out[6] VPWR VGND sg13g2_buf_1
XFILLER_0_203 VPWR VGND sg13g2_decap_8
XFILLER_29_410 VPWR VGND sg13g2_decap_8
XFILLER_45_936 VPWR VGND sg13g2_decap_8
XFILLER_17_616 VPWR VGND sg13g2_decap_8
XFILLER_29_487 VPWR VGND sg13g2_decap_8
XFILLER_44_446 VPWR VGND sg13g2_decap_8
XFILLER_16_137 VPWR VGND sg13g2_decap_8
XFILLER_13_844 VPWR VGND sg13g2_decap_8
XFILLER_12_354 VPWR VGND sg13g2_decap_8
XFILLER_40_663 VPWR VGND sg13g2_decap_8
XFILLER_9_837 VPWR VGND sg13g2_decap_8
XFILLER_8_347 VPWR VGND sg13g2_decap_8
XFILLER_21_81 VPWR VGND sg13g2_decap_8
XFILLER_4_564 VPWR VGND sg13g2_decap_8
XFILLER_39_207 VPWR VGND sg13g2_decap_8
XFILLER_0_770 VPWR VGND sg13g2_decap_8
XFILLER_48_763 VPWR VGND sg13g2_decap_8
XFILLER_47_273 VPWR VGND sg13g2_decap_8
XFILLER_35_402 VPWR VGND sg13g2_decap_8
XFILLER_36_914 VPWR VGND sg13g2_decap_8
XFILLER_35_479 VPWR VGND sg13g2_decap_8
XFILLER_16_671 VPWR VGND sg13g2_decap_8
XFILLER_31_652 VPWR VGND sg13g2_decap_8
XFILLER_30_173 VPWR VGND sg13g2_decap_8
XFILLER_11_1005 VPWR VGND sg13g2_decap_8
XFILLER_27_903 VPWR VGND sg13g2_decap_8
XFILLER_26_413 VPWR VGND sg13g2_decap_8
XFILLER_39_774 VPWR VGND sg13g2_decap_8
XFILLER_38_284 VPWR VGND sg13g2_decap_8
XFILLER_14_619 VPWR VGND sg13g2_decap_8
XFILLER_42_47 VPWR VGND sg13g2_decap_8
XFILLER_21_151 VPWR VGND sg13g2_decap_8
XFILLER_21_162 VPWR VGND sg13g2_decap_8
XFILLER_22_674 VPWR VGND sg13g2_decap_8
XFILLER_10_858 VPWR VGND sg13g2_decap_8
XFILLER_27_1001 VPWR VGND sg13g2_decap_8
XFILLER_1_567 VPWR VGND sg13g2_decap_8
XFILLER_17_413 VPWR VGND sg13g2_decap_8
XFILLER_18_914 VPWR VGND sg13g2_decap_8
XFILLER_45_733 VPWR VGND sg13g2_decap_8
XFILLER_44_243 VPWR VGND sg13g2_decap_8
XFILLER_26_980 VPWR VGND sg13g2_decap_8
XFILLER_41_950 VPWR VGND sg13g2_decap_8
XFILLER_13_641 VPWR VGND sg13g2_decap_8
XFILLER_16_81 VPWR VGND sg13g2_decap_8
XFILLER_9_634 VPWR VGND sg13g2_decap_8
XFILLER_12_151 VPWR VGND sg13g2_decap_8
XFILLER_40_460 VPWR VGND sg13g2_decap_8
XFILLER_8_144 VPWR VGND sg13g2_decap_8
XFILLER_5_851 VPWR VGND sg13g2_decap_8
XFILLER_4_361 VPWR VGND sg13g2_decap_8
XFILLER_48_560 VPWR VGND sg13g2_decap_8
XFILLER_36_711 VPWR VGND sg13g2_decap_8
XFILLER_35_221 VPWR VGND sg13g2_decap_8
XFILLER_24_928 VPWR VGND sg13g2_decap_8
XFILLER_36_788 VPWR VGND sg13g2_decap_8
XFILLER_17_980 VPWR VGND sg13g2_decap_8
XFILLER_23_438 VPWR VGND sg13g2_decap_8
XFILLER_32_950 VPWR VGND sg13g2_decap_8
XFILLER_12_39 VPWR VGND sg13g2_decap_8
XFILLER_37_14 VPWR VGND sg13g2_decap_8
XFILLER_27_700 VPWR VGND sg13g2_decap_8
XFILLER_39_571 VPWR VGND sg13g2_decap_8
XFILLER_26_221 VPWR VGND sg13g2_decap_8
XFILLER_15_917 VPWR VGND sg13g2_decap_8
XFILLER_27_777 VPWR VGND sg13g2_decap_8
XFILLER_42_747 VPWR VGND sg13g2_decap_8
XFILLER_14_416 VPWR VGND sg13g2_decap_8
XFILLER_41_235 VPWR VGND sg13g2_decap_8
XFILLER_22_471 VPWR VGND sg13g2_decap_8
XFILLER_10_655 VPWR VGND sg13g2_decap_8
XFILLER_6_648 VPWR VGND sg13g2_decap_8
XFILLER_5_158 VPWR VGND sg13g2_decap_8
XFILLER_2_865 VPWR VGND sg13g2_decap_8
XFILLER_1_364 VPWR VGND sg13g2_decap_8
XFILLER_49_357 VPWR VGND sg13g2_decap_8
XFILLER_18_711 VPWR VGND sg13g2_decap_8
XFILLER_40_1020 VPWR VGND sg13g2_decap_8
XFILLER_45_530 VPWR VGND sg13g2_decap_8
XFILLER_17_210 VPWR VGND sg13g2_decap_8
XFILLER_18_788 VPWR VGND sg13g2_decap_8
XFILLER_17_287 VPWR VGND sg13g2_decap_8
XFILLER_27_91 VPWR VGND sg13g2_decap_8
XFILLER_33_747 VPWR VGND sg13g2_decap_8
XFILLER_32_257 VPWR VGND sg13g2_decap_8
XFILLER_14_983 VPWR VGND sg13g2_decap_8
XFILLER_9_431 VPWR VGND sg13g2_decap_8
XFILLER_4_95 VPWR VGND sg13g2_decap_8
XFILLER_28_519 VPWR VGND sg13g2_decap_8
XFILLER_24_725 VPWR VGND sg13g2_decap_8
XFILLER_36_585 VPWR VGND sg13g2_decap_8
XFILLER_17_1022 VPWR VGND sg13g2_decap_8
XFILLER_20_964 VPWR VGND sg13g2_decap_8
XFILLER_48_35 VPWR VGND sg13g2_decap_8
XFILLER_24_1026 VPWR VGND sg13g2_fill_2
XFILLER_15_714 VPWR VGND sg13g2_decap_8
XFILLER_27_574 VPWR VGND sg13g2_decap_8
XFILLER_42_544 VPWR VGND sg13g2_decap_8
XFILLER_9_18 VPWR VGND sg13g2_decap_8
XFILLER_11_942 VPWR VGND sg13g2_decap_8
XFILLER_10_452 VPWR VGND sg13g2_decap_8
XFILLER_7_924 VPWR VGND sg13g2_decap_8
XFILLER_13_60 VPWR VGND sg13g2_decap_8
XFILLER_6_445 VPWR VGND sg13g2_decap_8
XFILLER_2_662 VPWR VGND sg13g2_decap_8
XFILLER_1_161 VPWR VGND sg13g2_decap_8
XFILLER_29_7 VPWR VGND sg13g2_decap_8
XFILLER_49_154 VPWR VGND sg13g2_decap_8
XFILLER_38_806 VPWR VGND sg13g2_decap_8
XFILLER_37_349 VPWR VGND sg13g2_decap_8
XFILLER_46_861 VPWR VGND sg13g2_decap_8
XFILLER_18_585 VPWR VGND sg13g2_decap_8
XFILLER_33_544 VPWR VGND sg13g2_decap_8
XFILLER_21_717 VPWR VGND sg13g2_decap_8
XFILLER_14_780 VPWR VGND sg13g2_decap_8
XFILLER_20_249 VPWR VGND sg13g2_decap_8
XFILLER_47_1015 VPWR VGND sg13g2_decap_8
XFILLER_24_522 VPWR VGND sg13g2_decap_8
XFILLER_34_26 VPWR VGND sg13g2_decap_8
XFILLER_36_382 VPWR VGND sg13g2_decap_8
XFILLER_12_739 VPWR VGND sg13g2_decap_8
XFILLER_24_599 VPWR VGND sg13g2_decap_8
XFILLER_11_249 VPWR VGND sg13g2_decap_8
XFILLER_20_761 VPWR VGND sg13g2_decap_8
XFILLER_4_949 VPWR VGND sg13g2_decap_8
XFILLER_3_459 VPWR VGND sg13g2_decap_8
XFILLER_47_658 VPWR VGND sg13g2_decap_8
XFILLER_46_168 VPWR VGND sg13g2_decap_8
XFILLER_15_511 VPWR VGND sg13g2_decap_8
XFILLER_27_371 VPWR VGND sg13g2_decap_8
XFILLER_28_883 VPWR VGND sg13g2_decap_8
XFILLER_43_831 VPWR VGND sg13g2_decap_8
XFILLER_42_341 VPWR VGND sg13g2_decap_8
XFILLER_15_588 VPWR VGND sg13g2_decap_8
XFILLER_24_81 VPWR VGND sg13g2_decap_8
XFILLER_30_569 VPWR VGND sg13g2_decap_8
XFILLER_7_721 VPWR VGND sg13g2_decap_8
XFILLER_6_242 VPWR VGND sg13g2_decap_8
XFILLER_7_798 VPWR VGND sg13g2_decap_8
X_098_ _020_ net3 net2 VPWR VGND sg13g2_nand2b_1
XFILLER_34_5 VPWR VGND sg13g2_decap_8
XFILLER_38_603 VPWR VGND sg13g2_decap_8
XFILLER_1_63 VPWR VGND sg13g2_decap_8
XFILLER_18_382 VPWR VGND sg13g2_decap_8
XFILLER_34_853 VPWR VGND sg13g2_decap_8
XFILLER_21_514 VPWR VGND sg13g2_decap_8
XFILLER_33_385 VPWR VGND sg13g2_decap_8
XFILLER_14_1025 VPWR VGND sg13g2_decap_4
XFILLER_20_39 VPWR VGND sg13g2_decap_8
XFILLER_21_1018 VPWR VGND sg13g2_decap_8
XFILLER_28_102 VPWR VGND sg13g2_decap_8
XFILLER_29_669 VPWR VGND sg13g2_decap_8
XFILLER_45_47 VPWR VGND sg13g2_decap_8
XFILLER_44_628 VPWR VGND sg13g2_decap_8
XFILLER_16_319 VPWR VGND sg13g2_decap_8
XFILLER_43_138 VPWR VGND sg13g2_decap_8
XFILLER_25_831 VPWR VGND sg13g2_decap_8
XFILLER_12_536 VPWR VGND sg13g2_decap_8
XFILLER_40_845 VPWR VGND sg13g2_decap_8
XFILLER_8_529 VPWR VGND sg13g2_decap_8
XFILLER_4_746 VPWR VGND sg13g2_decap_8
XFILLER_3_256 VPWR VGND sg13g2_decap_8
XFILLER_0_952 VPWR VGND sg13g2_decap_8
XFILLER_48_945 VPWR VGND sg13g2_decap_8
XFILLER_19_102 VPWR VGND sg13g2_decap_8
XFILLER_47_455 VPWR VGND sg13g2_decap_8
XFILLER_19_81 VPWR VGND sg13g2_decap_8
XFILLER_16_853 VPWR VGND sg13g2_decap_8
XFILLER_28_680 VPWR VGND sg13g2_decap_8
XFILLER_34_138 VPWR VGND sg13g2_decap_8
XFILLER_37_1014 VPWR VGND sg13g2_decap_8
XFILLER_15_385 VPWR VGND sg13g2_decap_8
XFILLER_30_311 VPWR VGND sg13g2_decap_8
XFILLER_31_834 VPWR VGND sg13g2_decap_8
XFILLER_30_366 VPWR VGND sg13g2_decap_8
XFILLER_7_595 VPWR VGND sg13g2_decap_8
Xheichips25_template_28 VPWR VGND uio_out[4] sg13g2_tielo
XFILLER_38_400 VPWR VGND sg13g2_decap_8
Xheichips25_template_39 VPWR VGND uio_oe[6] sg13g2_tiehi
XFILLER_39_956 VPWR VGND sg13g2_decap_8
XFILLER_38_477 VPWR VGND sg13g2_decap_8
XFILLER_25_116 VPWR VGND sg13g2_decap_8
XFILLER_15_39 VPWR VGND sg13g2_decap_8
XFILLER_34_650 VPWR VGND sg13g2_decap_8
XFILLER_22_856 VPWR VGND sg13g2_decap_8
XFILLER_33_182 VPWR VGND sg13g2_decap_8
XFILLER_21_388 VPWR VGND sg13g2_decap_8
Xoutput27 net32 uo_out[7] VPWR VGND sg13g2_buf_1
Xoutput16 net21 uio_out[0] VPWR VGND sg13g2_buf_1
XFILLER_1_749 VPWR VGND sg13g2_decap_8
XFILLER_0_259 VPWR VGND sg13g2_decap_8
XFILLER_5_1012 VPWR VGND sg13g2_decap_8
XFILLER_45_915 VPWR VGND sg13g2_decap_8
XFILLER_29_466 VPWR VGND sg13g2_decap_8
XFILLER_44_425 VPWR VGND sg13g2_decap_8
XFILLER_16_116 VPWR VGND sg13g2_decap_8
XFILLER_13_823 VPWR VGND sg13g2_decap_8
XFILLER_9_816 VPWR VGND sg13g2_decap_8
XFILLER_12_333 VPWR VGND sg13g2_decap_8
XFILLER_40_642 VPWR VGND sg13g2_decap_8
XFILLER_8_326 VPWR VGND sg13g2_decap_8
XFILLER_4_543 VPWR VGND sg13g2_decap_8
XFILLER_21_60 VPWR VGND sg13g2_decap_8
XFILLER_48_742 VPWR VGND sg13g2_decap_8
XFILLER_47_252 VPWR VGND sg13g2_decap_8
XFILLER_16_650 VPWR VGND sg13g2_decap_8
XFILLER_35_458 VPWR VGND sg13g2_decap_8
XFILLER_44_992 VPWR VGND sg13g2_decap_8
Xclkbuf_0_clk clk clknet_0_clk VPWR VGND sg13g2_buf_8
XFILLER_31_631 VPWR VGND sg13g2_decap_8
XFILLER_30_152 VPWR VGND sg13g2_decap_8
XFILLER_11_1028 VPWR VGND sg13g2_fill_1
XFILLER_8_893 VPWR VGND sg13g2_decap_8
XFILLER_7_392 VPWR VGND sg13g2_decap_8
XFILLER_7_84 VPWR VGND sg13g2_decap_8
XFILLER_39_753 VPWR VGND sg13g2_decap_8
XFILLER_38_263 VPWR VGND sg13g2_decap_8
XFILLER_27_959 VPWR VGND sg13g2_decap_8
XFILLER_42_929 VPWR VGND sg13g2_decap_8
XFILLER_26_469 VPWR VGND sg13g2_decap_8
XFILLER_41_439 VPWR VGND sg13g2_decap_8
XFILLER_42_26 VPWR VGND sg13g2_decap_8
XFILLER_21_130 VPWR VGND sg13g2_decap_8
XFILLER_22_653 VPWR VGND sg13g2_decap_8
XFILLER_10_837 VPWR VGND sg13g2_decap_8
XFILLER_1_546 VPWR VGND sg13g2_decap_8
XFILLER_49_539 VPWR VGND sg13g2_decap_8
XFILLER_45_712 VPWR VGND sg13g2_decap_8
XFILLER_44_222 VPWR VGND sg13g2_decap_8
XFILLER_29_285 VPWR VGND sg13g2_decap_4
XFILLER_29_296 VPWR VGND sg13g2_decap_8
XFILLER_45_789 VPWR VGND sg13g2_decap_8
XFILLER_17_469 VPWR VGND sg13g2_decap_8
XFILLER_33_929 VPWR VGND sg13g2_decap_8
XFILLER_44_299 VPWR VGND sg13g2_decap_8
XFILLER_16_60 VPWR VGND sg13g2_decap_8
XFILLER_32_439 VPWR VGND sg13g2_decap_8
XFILLER_13_620 VPWR VGND sg13g2_decap_8
XFILLER_9_613 VPWR VGND sg13g2_decap_8
XFILLER_12_130 VPWR VGND sg13g2_decap_8
XFILLER_34_1028 VPWR VGND sg13g2_fill_1
XFILLER_8_123 VPWR VGND sg13g2_decap_8
XFILLER_13_697 VPWR VGND sg13g2_decap_8
XFILLER_5_830 VPWR VGND sg13g2_decap_8
XFILLER_4_340 VPWR VGND sg13g2_decap_8
XFILLER_24_907 VPWR VGND sg13g2_decap_8
XFILLER_35_255 VPWR VGND sg13g2_decap_8
XFILLER_36_767 VPWR VGND sg13g2_decap_8
XFILLER_23_417 VPWR VGND sg13g2_decap_8
XFILLER_35_266 VPWR VGND sg13g2_fill_2
XFILLER_12_18 VPWR VGND sg13g2_decap_8
XFILLER_8_690 VPWR VGND sg13g2_decap_8
XFILLER_39_550 VPWR VGND sg13g2_decap_8
XFILLER_2_1026 VPWR VGND sg13g2_fill_2
XFILLER_26_200 VPWR VGND sg13g2_decap_8
XFILLER_27_756 VPWR VGND sg13g2_decap_8
XFILLER_42_726 VPWR VGND sg13g2_decap_8
XFILLER_26_288 VPWR VGND sg13g2_decap_8
XFILLER_41_214 VPWR VGND sg13g2_decap_8
XFILLER_22_450 VPWR VGND sg13g2_decap_8
XFILLER_23_984 VPWR VGND sg13g2_decap_8
XFILLER_10_634 VPWR VGND sg13g2_decap_8
XFILLER_6_627 VPWR VGND sg13g2_decap_8
XFILLER_5_137 VPWR VGND sg13g2_decap_8
XFILLER_2_844 VPWR VGND sg13g2_decap_8
XFILLER_1_343 VPWR VGND sg13g2_decap_8
XFILLER_49_336 VPWR VGND sg13g2_decap_8
XFILLER_18_767 VPWR VGND sg13g2_decap_8
XFILLER_27_70 VPWR VGND sg13g2_decap_8
XFILLER_45_586 VPWR VGND sg13g2_decap_8
XFILLER_17_266 VPWR VGND sg13g2_decap_8
XFILLER_33_726 VPWR VGND sg13g2_decap_8
XFILLER_32_236 VPWR VGND sg13g2_decap_8
XFILLER_9_410 VPWR VGND sg13g2_decap_8
XFILLER_14_962 VPWR VGND sg13g2_decap_8
XFILLER_13_494 VPWR VGND sg13g2_decap_8
XFILLER_9_487 VPWR VGND sg13g2_decap_8
XFILLER_4_74 VPWR VGND sg13g2_decap_8
XFILLER_24_704 VPWR VGND sg13g2_decap_8
XFILLER_36_564 VPWR VGND sg13g2_decap_8
XFILLER_17_1001 VPWR VGND sg13g2_decap_8
XFILLER_23_258 VPWR VGND sg13g2_decap_8
XFILLER_20_943 VPWR VGND sg13g2_decap_8
XFILLER_23_39 VPWR VGND sg13g2_decap_8
XFILLER_48_14 VPWR VGND sg13g2_decap_8
XFILLER_24_1005 VPWR VGND sg13g2_decap_8
XFILLER_27_553 VPWR VGND sg13g2_decap_8
XFILLER_42_523 VPWR VGND sg13g2_decap_8
XFILLER_14_214 VPWR VGND sg13g2_decap_8
XFILLER_14_269 VPWR VGND sg13g2_decap_8
XFILLER_11_921 VPWR VGND sg13g2_decap_8
XFILLER_23_781 VPWR VGND sg13g2_decap_8
XFILLER_10_431 VPWR VGND sg13g2_decap_8
XFILLER_7_903 VPWR VGND sg13g2_decap_8
XFILLER_31_1009 VPWR VGND sg13g2_decap_8
XFILLER_6_424 VPWR VGND sg13g2_decap_8
XFILLER_11_998 VPWR VGND sg13g2_decap_8
XFILLER_2_641 VPWR VGND sg13g2_decap_8
XFILLER_1_140 VPWR VGND sg13g2_decap_8
XFILLER_49_133 VPWR VGND sg13g2_decap_8
XFILLER_37_306 VPWR VGND sg13g2_decap_8
XFILLER_37_317 VPWR VGND sg13g2_fill_1
XFILLER_37_328 VPWR VGND sg13g2_decap_8
XFILLER_46_840 VPWR VGND sg13g2_decap_8
XFILLER_18_564 VPWR VGND sg13g2_decap_8
XFILLER_45_383 VPWR VGND sg13g2_decap_8
XFILLER_33_523 VPWR VGND sg13g2_decap_8
XFILLER_20_228 VPWR VGND sg13g2_decap_8
XFILLER_13_291 VPWR VGND sg13g2_decap_8
XFILLER_9_284 VPWR VGND sg13g2_decap_8
XFILLER_6_991 VPWR VGND sg13g2_decap_8
XFILLER_48_0 VPWR VGND sg13g2_decap_8
XFILLER_18_39 VPWR VGND sg13g2_decap_8
XFILLER_28_328 VPWR VGND sg13g2_fill_2
XFILLER_24_501 VPWR VGND sg13g2_decap_8
XFILLER_36_361 VPWR VGND sg13g2_decap_8
XFILLER_37_895 VPWR VGND sg13g2_decap_8
XFILLER_12_718 VPWR VGND sg13g2_decap_8
XFILLER_24_578 VPWR VGND sg13g2_decap_8
XFILLER_11_228 VPWR VGND sg13g2_decap_8
XFILLER_20_740 VPWR VGND sg13g2_decap_8
XFILLER_4_928 VPWR VGND sg13g2_decap_8
XFILLER_3_438 VPWR VGND sg13g2_decap_8
XFILLER_47_637 VPWR VGND sg13g2_decap_8
XFILLER_19_339 VPWR VGND sg13g2_decap_8
XFILLER_46_147 VPWR VGND sg13g2_decap_8
XFILLER_43_810 VPWR VGND sg13g2_decap_8
XFILLER_27_350 VPWR VGND sg13g2_decap_8
XFILLER_28_862 VPWR VGND sg13g2_decap_8
XFILLER_42_320 VPWR VGND sg13g2_decap_8
XFILLER_43_887 VPWR VGND sg13g2_decap_8
XFILLER_15_567 VPWR VGND sg13g2_decap_8
XFILLER_42_397 VPWR VGND sg13g2_decap_8
XFILLER_24_60 VPWR VGND sg13g2_decap_8
XFILLER_7_700 VPWR VGND sg13g2_decap_8
XFILLER_30_548 VPWR VGND sg13g2_decap_8
XFILLER_7_777 VPWR VGND sg13g2_decap_8
XFILLER_6_221 VPWR VGND sg13g2_decap_8
XFILLER_11_795 VPWR VGND sg13g2_decap_8
X_097_ mod1.qam16_mod.q_level\[3\] net2 _019_ VPWR VGND sg13g2_nor2_1
XFILLER_40_81 VPWR VGND sg13g2_decap_8
XFILLER_6_298 VPWR VGND sg13g2_decap_8
XFILLER_1_42 VPWR VGND sg13g2_decap_8
XFILLER_37_147 VPWR VGND sg13g2_decap_4
XFILLER_38_659 VPWR VGND sg13g2_decap_8
XFILLER_18_361 VPWR VGND sg13g2_decap_8
XFILLER_45_180 VPWR VGND sg13g2_decap_8
XFILLER_19_895 VPWR VGND sg13g2_decap_8
XFILLER_34_832 VPWR VGND sg13g2_decap_8
XFILLER_33_364 VPWR VGND sg13g2_decap_8
XFILLER_14_1004 VPWR VGND sg13g2_decap_8
XFILLER_20_18 VPWR VGND sg13g2_decap_8
XFILLER_29_49 VPWR VGND sg13g2_decap_8
XFILLER_29_648 VPWR VGND sg13g2_decap_8
XFILLER_45_26 VPWR VGND sg13g2_decap_8
XFILLER_44_607 VPWR VGND sg13g2_decap_8
XFILLER_25_810 VPWR VGND sg13g2_decap_8
XFILLER_43_117 VPWR VGND sg13g2_decap_8
XFILLER_24_320 VPWR VGND sg13g2_decap_8
XFILLER_36_180 VPWR VGND sg13g2_decap_8
XFILLER_37_692 VPWR VGND sg13g2_decap_8
XFILLER_25_887 VPWR VGND sg13g2_decap_8
XFILLER_12_515 VPWR VGND sg13g2_decap_8
XFILLER_24_386 VPWR VGND sg13g2_decap_8
XFILLER_40_824 VPWR VGND sg13g2_decap_8
XFILLER_8_508 VPWR VGND sg13g2_decap_8
XFILLER_4_725 VPWR VGND sg13g2_decap_8
XFILLER_3_235 VPWR VGND sg13g2_decap_8
XFILLER_10_95 VPWR VGND sg13g2_decap_8
XFILLER_0_931 VPWR VGND sg13g2_decap_8
XFILLER_48_924 VPWR VGND sg13g2_decap_8
XFILLER_47_434 VPWR VGND sg13g2_decap_8
XFILLER_19_60 VPWR VGND sg13g2_decap_8
XFILLER_16_832 VPWR VGND sg13g2_decap_8
XFILLER_34_117 VPWR VGND sg13g2_decap_8
XFILLER_43_684 VPWR VGND sg13g2_decap_8
XFILLER_15_364 VPWR VGND sg13g2_decap_8
XFILLER_31_813 VPWR VGND sg13g2_decap_8
XFILLER_42_194 VPWR VGND sg13g2_decap_8
XFILLER_30_334 VPWR VGND sg13g2_fill_1
XFILLER_11_592 VPWR VGND sg13g2_decap_8
XFILLER_7_574 VPWR VGND sg13g2_decap_8
XFILLER_39_935 VPWR VGND sg13g2_decap_8
Xheichips25_template_29 VPWR VGND uio_out[5] sg13g2_tielo
XFILLER_38_456 VPWR VGND sg13g2_decap_8
XFILLER_19_692 VPWR VGND sg13g2_decap_8
XFILLER_15_18 VPWR VGND sg13g2_decap_8
XFILLER_21_312 VPWR VGND sg13g2_decap_8
XFILLER_22_835 VPWR VGND sg13g2_decap_8
XFILLER_40_109 VPWR VGND sg13g2_decap_8
XFILLER_21_367 VPWR VGND sg13g2_decap_8
Xoutput17 net22 uio_out[1] VPWR VGND sg13g2_buf_1
XFILLER_1_728 VPWR VGND sg13g2_decap_8
XFILLER_0_238 VPWR VGND sg13g2_decap_8
XFILLER_29_445 VPWR VGND sg13g2_decap_8
XFILLER_44_404 VPWR VGND sg13g2_decap_8
XFILLER_13_802 VPWR VGND sg13g2_decap_8
XFILLER_12_312 VPWR VGND sg13g2_decap_8
XFILLER_24_172 VPWR VGND sg13g2_decap_8
XFILLER_25_684 VPWR VGND sg13g2_decap_8
XFILLER_40_621 VPWR VGND sg13g2_decap_8
XFILLER_8_305 VPWR VGND sg13g2_decap_8
XFILLER_13_879 VPWR VGND sg13g2_decap_8
XFILLER_12_389 VPWR VGND sg13g2_decap_8
XFILLER_40_698 VPWR VGND sg13g2_decap_8
XFILLER_4_522 VPWR VGND sg13g2_decap_8
XFILLER_4_599 VPWR VGND sg13g2_decap_8
XFILLER_48_721 VPWR VGND sg13g2_decap_8
XFILLER_47_231 VPWR VGND sg13g2_decap_8
XFILLER_48_798 VPWR VGND sg13g2_decap_8
XFILLER_35_437 VPWR VGND sg13g2_decap_8
XFILLER_36_949 VPWR VGND sg13g2_decap_8
XFILLER_46_91 VPWR VGND sg13g2_decap_8
XFILLER_44_971 VPWR VGND sg13g2_decap_8
XFILLER_22_109 VPWR VGND sg13g2_decap_8
XFILLER_31_610 VPWR VGND sg13g2_decap_8
XFILLER_43_481 VPWR VGND sg13g2_decap_8
XFILLER_15_172 VPWR VGND sg13g2_decap_4
XFILLER_30_131 VPWR VGND sg13g2_decap_8
XFILLER_31_687 VPWR VGND sg13g2_decap_8
XFILLER_8_872 VPWR VGND sg13g2_decap_8
XFILLER_7_63 VPWR VGND sg13g2_decap_8
XFILLER_7_371 VPWR VGND sg13g2_decap_8
XFILLER_39_732 VPWR VGND sg13g2_decap_8
XFILLER_38_242 VPWR VGND sg13g2_decap_8
XFILLER_26_39 VPWR VGND sg13g2_decap_8
XFILLER_27_938 VPWR VGND sg13g2_decap_8
XFILLER_42_908 VPWR VGND sg13g2_decap_8
XFILLER_26_448 VPWR VGND sg13g2_decap_8
XFILLER_41_418 VPWR VGND sg13g2_decap_8
XFILLER_13_109 VPWR VGND sg13g2_decap_8
XFILLER_22_632 VPWR VGND sg13g2_decap_8
XFILLER_10_816 VPWR VGND sg13g2_decap_8
XFILLER_6_809 VPWR VGND sg13g2_decap_8
XFILLER_21_197 VPWR VGND sg13g2_decap_8
XFILLER_5_319 VPWR VGND sg13g2_decap_8
XFILLER_1_525 VPWR VGND sg13g2_decap_8
XFILLER_49_518 VPWR VGND sg13g2_decap_8
XFILLER_29_264 VPWR VGND sg13g2_decap_8
XFILLER_44_201 VPWR VGND sg13g2_decap_8
XFILLER_18_949 VPWR VGND sg13g2_decap_8
XFILLER_45_768 VPWR VGND sg13g2_decap_8
XFILLER_17_448 VPWR VGND sg13g2_decap_8
XFILLER_33_908 VPWR VGND sg13g2_decap_8
XFILLER_44_278 VPWR VGND sg13g2_decap_8
XFILLER_32_418 VPWR VGND sg13g2_decap_8
XFILLER_25_481 VPWR VGND sg13g2_decap_8
XFILLER_41_985 VPWR VGND sg13g2_decap_8
XFILLER_8_102 VPWR VGND sg13g2_decap_8
XFILLER_13_676 VPWR VGND sg13g2_decap_8
XFILLER_34_1007 VPWR VGND sg13g2_decap_8
XFILLER_9_669 VPWR VGND sg13g2_decap_8
XFILLER_12_186 VPWR VGND sg13g2_decap_8
XFILLER_40_495 VPWR VGND sg13g2_decap_8
XFILLER_8_179 VPWR VGND sg13g2_decap_8
XFILLER_32_82 VPWR VGND sg13g2_decap_8
XFILLER_5_886 VPWR VGND sg13g2_decap_8
XFILLER_4_396 VPWR VGND sg13g2_decap_8
XFILLER_48_595 VPWR VGND sg13g2_decap_8
XFILLER_35_201 VPWR VGND sg13g2_fill_1
XFILLER_36_746 VPWR VGND sg13g2_decap_8
XFILLER_35_278 VPWR VGND sg13g2_decap_8
XFILLER_32_985 VPWR VGND sg13g2_decap_8
XFILLER_31_484 VPWR VGND sg13g2_decap_8
XFILLER_2_1005 VPWR VGND sg13g2_decap_8
XFILLER_37_49 VPWR VGND sg13g2_decap_8
XFILLER_27_735 VPWR VGND sg13g2_decap_8
XFILLER_42_705 VPWR VGND sg13g2_decap_8
XFILLER_26_267 VPWR VGND sg13g2_decap_8
XFILLER_23_963 VPWR VGND sg13g2_decap_8
XFILLER_10_613 VPWR VGND sg13g2_decap_8
XFILLER_6_606 VPWR VGND sg13g2_decap_8
XFILLER_5_116 VPWR VGND sg13g2_decap_8
XFILLER_2_823 VPWR VGND sg13g2_decap_8
XFILLER_1_322 VPWR VGND sg13g2_decap_8
XFILLER_49_315 VPWR VGND sg13g2_decap_8
XFILLER_1_399 VPWR VGND sg13g2_decap_8
XFILLER_17_245 VPWR VGND sg13g2_decap_8
XFILLER_18_746 VPWR VGND sg13g2_decap_8
XFILLER_45_565 VPWR VGND sg13g2_decap_8
Xclkbuf_2_0__f_clk clknet_0_clk clknet_2_0__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_33_705 VPWR VGND sg13g2_decap_8
XFILLER_14_941 VPWR VGND sg13g2_decap_8
XFILLER_32_215 VPWR VGND sg13g2_decap_8
XFILLER_41_782 VPWR VGND sg13g2_decap_8
XFILLER_13_473 VPWR VGND sg13g2_decap_8
XFILLER_9_466 VPWR VGND sg13g2_decap_8
XFILLER_5_683 VPWR VGND sg13g2_decap_8
XFILLER_4_193 VPWR VGND sg13g2_decap_8
XFILLER_4_53 VPWR VGND sg13g2_decap_8
XFILLER_49_882 VPWR VGND sg13g2_decap_8
XFILLER_48_392 VPWR VGND sg13g2_decap_8
XFILLER_36_543 VPWR VGND sg13g2_decap_8
XFILLER_23_204 VPWR VGND sg13g2_decap_8
XFILLER_23_237 VPWR VGND sg13g2_decap_8
XFILLER_23_18 VPWR VGND sg13g2_decap_8
XFILLER_20_922 VPWR VGND sg13g2_decap_8
XFILLER_32_782 VPWR VGND sg13g2_decap_8
XFILLER_31_281 VPWR VGND sg13g2_decap_8
XFILLER_20_999 VPWR VGND sg13g2_decap_8
XFILLER_47_819 VPWR VGND sg13g2_decap_8
XFILLER_24_1028 VPWR VGND sg13g2_fill_1
XFILLER_46_329 VPWR VGND sg13g2_decap_8
XFILLER_27_532 VPWR VGND sg13g2_decap_8
XFILLER_42_502 VPWR VGND sg13g2_decap_8
XFILLER_15_749 VPWR VGND sg13g2_decap_8
XFILLER_42_579 VPWR VGND sg13g2_decap_8
XFILLER_11_900 VPWR VGND sg13g2_decap_8
XFILLER_23_760 VPWR VGND sg13g2_decap_8
XFILLER_10_410 VPWR VGND sg13g2_decap_8
XFILLER_11_977 VPWR VGND sg13g2_decap_8
XFILLER_10_487 VPWR VGND sg13g2_decap_8
XFILLER_7_959 VPWR VGND sg13g2_decap_8
XFILLER_6_403 VPWR VGND sg13g2_decap_8
XFILLER_13_95 VPWR VGND sg13g2_decap_8
XFILLER_2_620 VPWR VGND sg13g2_decap_8
XFILLER_49_112 VPWR VGND sg13g2_decap_8
XFILLER_2_697 VPWR VGND sg13g2_decap_8
XFILLER_1_196 VPWR VGND sg13g2_decap_8
XFILLER_49_189 VPWR VGND sg13g2_decap_8
XFILLER_38_81 VPWR VGND sg13g2_decap_8
XFILLER_18_543 VPWR VGND sg13g2_decap_8
XFILLER_46_896 VPWR VGND sg13g2_decap_8
XFILLER_45_362 VPWR VGND sg13g2_decap_8
XFILLER_33_502 VPWR VGND sg13g2_decap_8
XFILLER_33_579 VPWR VGND sg13g2_decap_8
XFILLER_13_270 VPWR VGND sg13g2_decap_8
XFILLER_20_207 VPWR VGND sg13g2_decap_8
XFILLER_9_263 VPWR VGND sg13g2_decap_8
XFILLER_6_970 VPWR VGND sg13g2_decap_8
XFILLER_5_480 VPWR VGND sg13g2_decap_8
XFILLER_18_18 VPWR VGND sg13g2_decap_8
XFILLER_28_307 VPWR VGND sg13g2_decap_8
XFILLER_36_340 VPWR VGND sg13g2_decap_8
XFILLER_37_874 VPWR VGND sg13g2_decap_8
XFILLER_24_557 VPWR VGND sg13g2_decap_8
XFILLER_11_207 VPWR VGND sg13g2_decap_8
XFILLER_30_1010 VPWR VGND sg13g2_decap_8
XFILLER_4_907 VPWR VGND sg13g2_decap_8
XFILLER_20_796 VPWR VGND sg13g2_decap_8
XFILLER_3_417 VPWR VGND sg13g2_decap_8
XFILLER_1_7 VPWR VGND sg13g2_decap_8
XFILLER_47_616 VPWR VGND sg13g2_decap_8
XFILLER_19_318 VPWR VGND sg13g2_decap_8
XFILLER_46_126 VPWR VGND sg13g2_decap_8
XFILLER_28_841 VPWR VGND sg13g2_decap_8
XFILLER_43_866 VPWR VGND sg13g2_decap_8
XFILLER_15_546 VPWR VGND sg13g2_decap_8
XFILLER_42_376 VPWR VGND sg13g2_decap_8
XFILLER_30_527 VPWR VGND sg13g2_decap_8
XFILLER_6_200 VPWR VGND sg13g2_decap_8
XFILLER_11_774 VPWR VGND sg13g2_decap_8
XFILLER_10_284 VPWR VGND sg13g2_decap_8
XFILLER_7_756 VPWR VGND sg13g2_decap_8
XFILLER_6_277 VPWR VGND sg13g2_decap_8
X_096_ net32 _016_ _018_ VPWR VGND sg13g2_nand2_2
XFILLER_40_60 VPWR VGND sg13g2_decap_8
XFILLER_3_984 VPWR VGND sg13g2_decap_8
XFILLER_49_91 VPWR VGND sg13g2_decap_8
XFILLER_2_494 VPWR VGND sg13g2_decap_8
XFILLER_1_21 VPWR VGND sg13g2_decap_8
XFILLER_38_638 VPWR VGND sg13g2_decap_8
XFILLER_37_126 VPWR VGND sg13g2_decap_8
XFILLER_1_98 VPWR VGND sg13g2_decap_8
XFILLER_18_340 VPWR VGND sg13g2_decap_8
XFILLER_19_874 VPWR VGND sg13g2_decap_8
XFILLER_34_811 VPWR VGND sg13g2_decap_8
XFILLER_46_693 VPWR VGND sg13g2_decap_8
XFILLER_34_888 VPWR VGND sg13g2_decap_8
XFILLER_21_549 VPWR VGND sg13g2_decap_8
XFILLER_29_28 VPWR VGND sg13g2_decap_8
XFILLER_29_627 VPWR VGND sg13g2_decap_8
XFILLER_28_137 VPWR VGND sg13g2_decap_8
XFILLER_28_148 VPWR VGND sg13g2_fill_1
XFILLER_37_671 VPWR VGND sg13g2_decap_8
XFILLER_25_866 VPWR VGND sg13g2_decap_8
XFILLER_40_803 VPWR VGND sg13g2_decap_8
XFILLER_24_365 VPWR VGND sg13g2_decap_8
XFILLER_20_593 VPWR VGND sg13g2_decap_8
XFILLER_4_704 VPWR VGND sg13g2_decap_8
XFILLER_3_214 VPWR VGND sg13g2_decap_8
XFILLER_10_74 VPWR VGND sg13g2_decap_8
XFILLER_0_910 VPWR VGND sg13g2_decap_8
XFILLER_48_903 VPWR VGND sg13g2_decap_8
XFILLER_47_413 VPWR VGND sg13g2_decap_8
XFILLER_0_987 VPWR VGND sg13g2_decap_8
XFILLER_19_137 VPWR VGND sg13g2_decap_8
XFILLER_35_619 VPWR VGND sg13g2_decap_8
XFILLER_16_811 VPWR VGND sg13g2_decap_8
XFILLER_43_663 VPWR VGND sg13g2_decap_8
XFILLER_15_343 VPWR VGND sg13g2_decap_8
XFILLER_42_173 VPWR VGND sg13g2_decap_8
XFILLER_16_888 VPWR VGND sg13g2_decap_8
XFILLER_35_82 VPWR VGND sg13g2_decap_8
XFILLER_31_869 VPWR VGND sg13g2_decap_8
XFILLER_11_571 VPWR VGND sg13g2_decap_8
XFILLER_7_553 VPWR VGND sg13g2_decap_8
X_079_ _046_ _045_ mod1.i_out_qpsk\[1\] net11 Demo1.qam16_bits\[3\] VPWR VGND sg13g2_a22oi_1
XFILLER_3_781 VPWR VGND sg13g2_decap_8
XFILLER_2_291 VPWR VGND sg13g2_decap_8
XFILLER_39_914 VPWR VGND sg13g2_decap_8
XFILLER_38_435 VPWR VGND sg13g2_decap_8
XFILLER_20_1020 VPWR VGND sg13g2_decap_8
XFILLER_47_980 VPWR VGND sg13g2_decap_8
XFILLER_19_671 VPWR VGND sg13g2_decap_8
XFILLER_46_490 VPWR VGND sg13g2_decap_8
XFILLER_22_814 VPWR VGND sg13g2_decap_8
XFILLER_34_685 VPWR VGND sg13g2_decap_8
XFILLER_30_891 VPWR VGND sg13g2_decap_8
XFILLER_1_707 VPWR VGND sg13g2_decap_8
Xoutput18 net23 uio_out[2] VPWR VGND sg13g2_buf_1
XFILLER_0_217 VPWR VGND sg13g2_decap_8
XFILLER_29_424 VPWR VGND sg13g2_decap_8
XFILLER_24_151 VPWR VGND sg13g2_decap_8
XFILLER_25_663 VPWR VGND sg13g2_decap_8
XFILLER_40_600 VPWR VGND sg13g2_decap_8
XFILLER_13_858 VPWR VGND sg13g2_decap_8
XFILLER_12_368 VPWR VGND sg13g2_decap_8
XFILLER_40_677 VPWR VGND sg13g2_decap_8
XFILLER_4_501 VPWR VGND sg13g2_decap_8
XFILLER_21_95 VPWR VGND sg13g2_decap_8
XFILLER_4_578 VPWR VGND sg13g2_decap_8
XFILLER_48_700 VPWR VGND sg13g2_decap_8
XFILLER_43_1020 VPWR VGND sg13g2_decap_8
XFILLER_47_210 VPWR VGND sg13g2_decap_8
XFILLER_0_784 VPWR VGND sg13g2_decap_8
XFILLER_48_777 VPWR VGND sg13g2_decap_8
XFILLER_36_928 VPWR VGND sg13g2_decap_8
XFILLER_47_287 VPWR VGND sg13g2_decap_8
XFILLER_46_70 VPWR VGND sg13g2_decap_8
XFILLER_29_991 VPWR VGND sg13g2_decap_8
XFILLER_35_416 VPWR VGND sg13g2_decap_8
XFILLER_44_950 VPWR VGND sg13g2_decap_8
XFILLER_43_460 VPWR VGND sg13g2_decap_8
XFILLER_15_151 VPWR VGND sg13g2_decap_8
XFILLER_16_685 VPWR VGND sg13g2_decap_8
XFILLER_30_110 VPWR VGND sg13g2_decap_8
XFILLER_31_666 VPWR VGND sg13g2_decap_8
XFILLER_30_187 VPWR VGND sg13g2_decap_8
XFILLER_8_851 VPWR VGND sg13g2_decap_8
XFILLER_7_350 VPWR VGND sg13g2_decap_8
XFILLER_7_42 VPWR VGND sg13g2_decap_8
XFILLER_11_1019 VPWR VGND sg13g2_decap_8
XFILLER_39_711 VPWR VGND sg13g2_decap_8
XFILLER_38_221 VPWR VGND sg13g2_decap_8
XFILLER_27_917 VPWR VGND sg13g2_decap_8
XFILLER_39_788 VPWR VGND sg13g2_decap_8
XFILLER_26_18 VPWR VGND sg13g2_decap_8
XFILLER_26_427 VPWR VGND sg13g2_decap_8
XFILLER_38_298 VPWR VGND sg13g2_decap_8
XFILLER_22_611 VPWR VGND sg13g2_decap_8
XFILLER_35_983 VPWR VGND sg13g2_decap_8
XFILLER_34_482 VPWR VGND sg13g2_decap_8
XFILLER_21_176 VPWR VGND sg13g2_decap_8
XFILLER_22_688 VPWR VGND sg13g2_decap_8
XFILLER_1_504 VPWR VGND sg13g2_decap_8
XFILLER_27_1015 VPWR VGND sg13g2_decap_8
XFILLER_29_243 VPWR VGND sg13g2_decap_8
XFILLER_17_427 VPWR VGND sg13g2_decap_8
XFILLER_18_928 VPWR VGND sg13g2_decap_8
XFILLER_45_747 VPWR VGND sg13g2_decap_8
XFILLER_44_257 VPWR VGND sg13g2_decap_8
XFILLER_25_460 VPWR VGND sg13g2_decap_8
XFILLER_26_994 VPWR VGND sg13g2_decap_8
XFILLER_16_95 VPWR VGND sg13g2_decap_8
XFILLER_41_964 VPWR VGND sg13g2_decap_8
XFILLER_13_655 VPWR VGND sg13g2_decap_8
XFILLER_9_648 VPWR VGND sg13g2_decap_8
XFILLER_12_165 VPWR VGND sg13g2_decap_8
XFILLER_40_474 VPWR VGND sg13g2_decap_8
XFILLER_8_158 VPWR VGND sg13g2_decap_8
XFILLER_32_61 VPWR VGND sg13g2_decap_8
XFILLER_5_865 VPWR VGND sg13g2_decap_8
XFILLER_4_375 VPWR VGND sg13g2_decap_8
XFILLER_0_581 VPWR VGND sg13g2_decap_8
XFILLER_48_574 VPWR VGND sg13g2_decap_8
XFILLER_36_725 VPWR VGND sg13g2_decap_8
XFILLER_35_235 VPWR VGND sg13g2_fill_1
XFILLER_16_482 VPWR VGND sg13g2_decap_8
XFILLER_17_994 VPWR VGND sg13g2_decap_8
XFILLER_32_964 VPWR VGND sg13g2_decap_8
XFILLER_31_463 VPWR VGND sg13g2_decap_8
XFILLER_37_28 VPWR VGND sg13g2_decap_8
XFILLER_2_1028 VPWR VGND sg13g2_fill_1
XFILLER_27_714 VPWR VGND sg13g2_decap_8
XFILLER_39_585 VPWR VGND sg13g2_decap_8
XFILLER_26_246 VPWR VGND sg13g2_decap_8
XFILLER_23_942 VPWR VGND sg13g2_decap_8
XFILLER_35_780 VPWR VGND sg13g2_decap_8
XFILLER_41_249 VPWR VGND sg13g2_decap_8
XFILLER_22_485 VPWR VGND sg13g2_decap_8
XFILLER_10_669 VPWR VGND sg13g2_decap_8
XFILLER_2_802 VPWR VGND sg13g2_decap_8
XFILLER_1_301 VPWR VGND sg13g2_decap_8
XFILLER_2_879 VPWR VGND sg13g2_decap_8
XFILLER_1_378 VPWR VGND sg13g2_decap_8
XFILLER_18_725 VPWR VGND sg13g2_decap_8
XFILLER_45_544 VPWR VGND sg13g2_decap_8
XFILLER_17_224 VPWR VGND sg13g2_decap_8
XFILLER_14_920 VPWR VGND sg13g2_decap_8
XFILLER_26_791 VPWR VGND sg13g2_decap_8
XFILLER_41_761 VPWR VGND sg13g2_decap_8
XFILLER_13_452 VPWR VGND sg13g2_decap_8
XFILLER_25_290 VPWR VGND sg13g2_decap_8
XFILLER_43_82 VPWR VGND sg13g2_decap_8
XFILLER_14_997 VPWR VGND sg13g2_decap_8
XFILLER_40_271 VPWR VGND sg13g2_fill_1
XFILLER_9_445 VPWR VGND sg13g2_decap_8
XFILLER_5_662 VPWR VGND sg13g2_decap_8
XFILLER_4_172 VPWR VGND sg13g2_decap_8
XFILLER_4_32 VPWR VGND sg13g2_decap_8
XFILLER_49_861 VPWR VGND sg13g2_decap_8
XFILLER_48_371 VPWR VGND sg13g2_decap_8
XFILLER_36_522 VPWR VGND sg13g2_decap_8
XFILLER_17_791 VPWR VGND sg13g2_decap_8
XFILLER_24_739 VPWR VGND sg13g2_decap_8
XFILLER_36_599 VPWR VGND sg13g2_decap_8
XFILLER_20_901 VPWR VGND sg13g2_decap_8
XFILLER_32_761 VPWR VGND sg13g2_decap_8
XFILLER_31_260 VPWR VGND sg13g2_decap_8
XFILLER_20_978 VPWR VGND sg13g2_decap_8
XFILLER_2_109 VPWR VGND sg13g2_decap_8
XFILLER_48_49 VPWR VGND sg13g2_decap_8
XFILLER_46_308 VPWR VGND sg13g2_decap_8
XFILLER_27_511 VPWR VGND sg13g2_decap_8
XFILLER_39_382 VPWR VGND sg13g2_decap_8
XFILLER_15_728 VPWR VGND sg13g2_decap_8
XFILLER_27_588 VPWR VGND sg13g2_decap_8
XFILLER_42_558 VPWR VGND sg13g2_decap_8
XFILLER_30_709 VPWR VGND sg13g2_decap_8
XFILLER_11_956 VPWR VGND sg13g2_decap_8
XFILLER_10_466 VPWR VGND sg13g2_decap_8
XFILLER_7_938 VPWR VGND sg13g2_decap_8
XFILLER_13_74 VPWR VGND sg13g2_decap_8
XFILLER_6_459 VPWR VGND sg13g2_decap_8
XFILLER_2_676 VPWR VGND sg13g2_decap_8
XFILLER_1_175 VPWR VGND sg13g2_decap_8
XFILLER_49_168 VPWR VGND sg13g2_decap_8
XFILLER_38_60 VPWR VGND sg13g2_decap_8
XFILLER_18_522 VPWR VGND sg13g2_decap_8
XFILLER_46_875 VPWR VGND sg13g2_decap_8
XFILLER_45_341 VPWR VGND sg13g2_decap_8
XFILLER_18_599 VPWR VGND sg13g2_decap_8
XFILLER_33_558 VPWR VGND sg13g2_decap_8
XFILLER_9_242 VPWR VGND sg13g2_decap_8
XFILLER_14_794 VPWR VGND sg13g2_decap_8
XFILLER_29_809 VPWR VGND sg13g2_decap_8
XFILLER_37_853 VPWR VGND sg13g2_decap_8
XFILLER_24_536 VPWR VGND sg13g2_decap_8
XFILLER_36_396 VPWR VGND sg13g2_decap_8
XFILLER_20_775 VPWR VGND sg13g2_decap_8
XFILLER_8_1012 VPWR VGND sg13g2_decap_8
XFILLER_46_105 VPWR VGND sg13g2_decap_8
XFILLER_28_820 VPWR VGND sg13g2_decap_8
XFILLER_43_845 VPWR VGND sg13g2_decap_8
XFILLER_15_525 VPWR VGND sg13g2_decap_8
XFILLER_27_385 VPWR VGND sg13g2_decap_8
XFILLER_28_897 VPWR VGND sg13g2_decap_8
XFILLER_42_355 VPWR VGND sg13g2_decap_8
XFILLER_30_506 VPWR VGND sg13g2_decap_8
XFILLER_11_753 VPWR VGND sg13g2_decap_8
XFILLER_24_95 VPWR VGND sg13g2_decap_8
XFILLER_10_263 VPWR VGND sg13g2_decap_8
XFILLER_7_735 VPWR VGND sg13g2_decap_8
XFILLER_6_256 VPWR VGND sg13g2_decap_8
X_095_ _018_ mod1.q_out_qam16\[3\] net11 VPWR VGND sg13g2_nand2_1
XFILLER_3_963 VPWR VGND sg13g2_decap_8
XFILLER_2_473 VPWR VGND sg13g2_decap_8
XFILLER_49_70 VPWR VGND sg13g2_decap_8
XFILLER_27_7 VPWR VGND sg13g2_decap_8
XFILLER_37_105 VPWR VGND sg13g2_decap_8
XFILLER_38_617 VPWR VGND sg13g2_decap_8
XFILLER_1_77 VPWR VGND sg13g2_decap_8
XFILLER_19_853 VPWR VGND sg13g2_decap_8
XFILLER_46_672 VPWR VGND sg13g2_decap_8
XFILLER_18_396 VPWR VGND sg13g2_decap_8
XFILLER_33_333 VPWR VGND sg13g2_decap_8
XFILLER_34_867 VPWR VGND sg13g2_decap_8
XFILLER_21_528 VPWR VGND sg13g2_decap_8
XFILLER_14_591 VPWR VGND sg13g2_decap_8
XFILLER_33_399 VPWR VGND sg13g2_decap_4
XFILLER_29_606 VPWR VGND sg13g2_decap_8
XFILLER_28_116 VPWR VGND sg13g2_decap_8
XFILLER_37_650 VPWR VGND sg13g2_decap_8
XFILLER_25_845 VPWR VGND sg13g2_decap_8
XFILLER_40_859 VPWR VGND sg13g2_decap_8
XFILLER_20_572 VPWR VGND sg13g2_decap_8
XFILLER_10_53 VPWR VGND sg13g2_decap_8
XFILLER_0_966 VPWR VGND sg13g2_decap_8
XFILLER_48_959 VPWR VGND sg13g2_decap_8
XFILLER_19_116 VPWR VGND sg13g2_decap_8
XFILLER_47_469 VPWR VGND sg13g2_decap_8
XFILLER_19_95 VPWR VGND sg13g2_decap_8
XFILLER_28_694 VPWR VGND sg13g2_decap_8
XFILLER_43_642 VPWR VGND sg13g2_decap_8
XFILLER_16_867 VPWR VGND sg13g2_decap_8
XFILLER_27_182 VPWR VGND sg13g2_decap_8
XFILLER_35_61 VPWR VGND sg13g2_decap_8
XFILLER_42_152 VPWR VGND sg13g2_decap_8
XFILLER_37_1028 VPWR VGND sg13g2_fill_1
XFILLER_15_399 VPWR VGND sg13g2_decap_8
XFILLER_30_325 VPWR VGND sg13g2_decap_8
XFILLER_31_848 VPWR VGND sg13g2_decap_8
XFILLER_11_550 VPWR VGND sg13g2_decap_8
XFILLER_7_532 VPWR VGND sg13g2_decap_8
X_078_ net7 net6 _045_ VPWR VGND sg13g2_nor2b_2
XFILLER_3_760 VPWR VGND sg13g2_decap_8
XFILLER_2_270 VPWR VGND sg13g2_decap_8
XFILLER_32_5 VPWR VGND sg13g2_decap_8
XFILLER_25_4 VPWR VGND sg13g2_decap_8
XFILLER_38_414 VPWR VGND sg13g2_decap_8
XFILLER_19_650 VPWR VGND sg13g2_decap_8
XFILLER_26_609 VPWR VGND sg13g2_decap_8
XFILLER_18_193 VPWR VGND sg13g2_decap_8
XFILLER_34_664 VPWR VGND sg13g2_decap_8
XFILLER_33_196 VPWR VGND sg13g2_decap_8
XFILLER_30_870 VPWR VGND sg13g2_decap_8
XFILLER_31_19 VPWR VGND sg13g2_decap_8
Xoutput19 net24 uio_out[3] VPWR VGND sg13g2_buf_1
XFILLER_29_403 VPWR VGND sg13g2_decap_8
XFILLER_5_1026 VPWR VGND sg13g2_fill_2
XFILLER_45_929 VPWR VGND sg13g2_decap_8
XFILLER_17_609 VPWR VGND sg13g2_decap_8
XFILLER_44_439 VPWR VGND sg13g2_decap_8
XFILLER_38_981 VPWR VGND sg13g2_decap_8
XFILLER_25_642 VPWR VGND sg13g2_decap_8
XFILLER_24_130 VPWR VGND sg13g2_decap_8
XFILLER_13_837 VPWR VGND sg13g2_decap_8
XFILLER_12_347 VPWR VGND sg13g2_decap_8
XFILLER_40_656 VPWR VGND sg13g2_decap_8
XFILLER_21_892 VPWR VGND sg13g2_decap_8
XFILLER_20_391 VPWR VGND sg13g2_decap_4
XFILLER_4_557 VPWR VGND sg13g2_decap_8
XFILLER_21_74 VPWR VGND sg13g2_decap_8
XFILLER_0_763 VPWR VGND sg13g2_decap_8
XFILLER_48_756 VPWR VGND sg13g2_decap_8
XFILLER_36_907 VPWR VGND sg13g2_decap_8
XFILLER_47_266 VPWR VGND sg13g2_decap_8
XFILLER_29_970 VPWR VGND sg13g2_decap_8
XFILLER_28_491 VPWR VGND sg13g2_decap_8
XFILLER_15_130 VPWR VGND sg13g2_decap_8
XFILLER_16_664 VPWR VGND sg13g2_decap_8
XFILLER_31_645 VPWR VGND sg13g2_decap_8
XFILLER_8_830 VPWR VGND sg13g2_decap_8
XFILLER_7_21 VPWR VGND sg13g2_decap_8
XFILLER_30_166 VPWR VGND sg13g2_decap_8
XFILLER_7_98 VPWR VGND sg13g2_decap_8
XFILLER_38_200 VPWR VGND sg13g2_decap_8
XFILLER_39_767 VPWR VGND sg13g2_decap_8
XFILLER_26_406 VPWR VGND sg13g2_decap_8
XFILLER_38_277 VPWR VGND sg13g2_decap_8
XFILLER_34_461 VPWR VGND sg13g2_decap_8
XFILLER_35_962 VPWR VGND sg13g2_decap_8
XFILLER_21_144 VPWR VGND sg13g2_decap_8
XFILLER_22_667 VPWR VGND sg13g2_decap_8
XFILLER_18_907 VPWR VGND sg13g2_decap_8
XFILLER_29_222 VPWR VGND sg13g2_decap_8
XFILLER_45_726 VPWR VGND sg13g2_decap_8
XFILLER_17_406 VPWR VGND sg13g2_decap_8
XFILLER_44_236 VPWR VGND sg13g2_decap_8
XFILLER_26_973 VPWR VGND sg13g2_decap_8
XFILLER_41_943 VPWR VGND sg13g2_decap_8
XFILLER_13_634 VPWR VGND sg13g2_decap_8
XFILLER_16_74 VPWR VGND sg13g2_decap_8
XFILLER_12_144 VPWR VGND sg13g2_decap_8
XFILLER_40_453 VPWR VGND sg13g2_decap_8
XFILLER_9_627 VPWR VGND sg13g2_decap_8
XFILLER_32_40 VPWR VGND sg13g2_decap_8
XFILLER_8_137 VPWR VGND sg13g2_decap_8
XFILLER_5_844 VPWR VGND sg13g2_decap_8
XFILLER_4_354 VPWR VGND sg13g2_decap_8
XFILLER_0_560 VPWR VGND sg13g2_decap_8
XFILLER_48_553 VPWR VGND sg13g2_decap_8
XFILLER_36_704 VPWR VGND sg13g2_decap_8
XFILLER_35_214 VPWR VGND sg13g2_decap_8
XFILLER_17_973 VPWR VGND sg13g2_decap_8
XFILLER_16_461 VPWR VGND sg13g2_decap_8
XFILLER_32_943 VPWR VGND sg13g2_decap_8
XFILLER_31_442 VPWR VGND sg13g2_decap_8
XFILLER_39_564 VPWR VGND sg13g2_decap_8
XFILLER_26_214 VPWR VGND sg13g2_decap_8
XFILLER_14_409 VPWR VGND sg13g2_decap_8
XFILLER_23_921 VPWR VGND sg13g2_decap_8
XFILLER_41_228 VPWR VGND sg13g2_decap_8
XFILLER_34_280 VPWR VGND sg13g2_decap_8
XFILLER_22_464 VPWR VGND sg13g2_decap_8
XFILLER_23_998 VPWR VGND sg13g2_decap_8
XFILLER_33_1020 VPWR VGND sg13g2_decap_8
XFILLER_10_648 VPWR VGND sg13g2_decap_8
XFILLER_2_858 VPWR VGND sg13g2_decap_8
XFILLER_1_357 VPWR VGND sg13g2_decap_8
XFILLER_40_1013 VPWR VGND sg13g2_decap_8
XFILLER_17_203 VPWR VGND sg13g2_decap_8
XFILLER_18_704 VPWR VGND sg13g2_decap_8
XFILLER_45_523 VPWR VGND sg13g2_decap_8
XFILLER_27_84 VPWR VGND sg13g2_decap_8
XFILLER_26_770 VPWR VGND sg13g2_decap_8
XFILLER_41_740 VPWR VGND sg13g2_decap_8
XFILLER_13_431 VPWR VGND sg13g2_decap_8
XFILLER_14_976 VPWR VGND sg13g2_decap_8
XFILLER_43_61 VPWR VGND sg13g2_decap_8
XFILLER_9_424 VPWR VGND sg13g2_decap_8
XFILLER_40_250 VPWR VGND sg13g2_decap_8
XFILLER_5_641 VPWR VGND sg13g2_decap_8
XFILLER_4_151 VPWR VGND sg13g2_decap_8
XFILLER_4_11 VPWR VGND sg13g2_decap_8
XFILLER_4_88 VPWR VGND sg13g2_decap_8
XFILLER_49_840 VPWR VGND sg13g2_decap_8
XFILLER_48_350 VPWR VGND sg13g2_decap_8
XFILLER_36_501 VPWR VGND sg13g2_decap_8
XFILLER_24_718 VPWR VGND sg13g2_decap_8
XFILLER_36_578 VPWR VGND sg13g2_decap_8
XFILLER_17_770 VPWR VGND sg13g2_decap_8
XFILLER_16_291 VPWR VGND sg13g2_decap_8
XFILLER_17_1015 VPWR VGND sg13g2_decap_8
XFILLER_32_740 VPWR VGND sg13g2_decap_8
XFILLER_20_957 VPWR VGND sg13g2_decap_8
XFILLER_9_991 VPWR VGND sg13g2_decap_8
XFILLER_48_28 VPWR VGND sg13g2_decap_8
XFILLER_24_1019 VPWR VGND sg13g2_decap_8
XFILLER_39_361 VPWR VGND sg13g2_decap_8
XFILLER_15_707 VPWR VGND sg13g2_decap_8
XFILLER_27_567 VPWR VGND sg13g2_decap_8
XFILLER_42_537 VPWR VGND sg13g2_decap_8
XFILLER_22_261 VPWR VGND sg13g2_decap_8
XFILLER_7_917 VPWR VGND sg13g2_decap_8
XFILLER_11_935 VPWR VGND sg13g2_decap_8
XFILLER_23_795 VPWR VGND sg13g2_decap_8
XFILLER_10_445 VPWR VGND sg13g2_decap_8
XFILLER_13_53 VPWR VGND sg13g2_decap_8
XFILLER_6_438 VPWR VGND sg13g2_decap_8
XFILLER_2_655 VPWR VGND sg13g2_decap_8
XFILLER_1_154 VPWR VGND sg13g2_decap_8
XFILLER_49_147 VPWR VGND sg13g2_decap_8
XFILLER_18_501 VPWR VGND sg13g2_decap_8
XFILLER_45_320 VPWR VGND sg13g2_decap_8
XFILLER_46_854 VPWR VGND sg13g2_decap_8
XFILLER_18_578 VPWR VGND sg13g2_decap_8
XFILLER_45_397 VPWR VGND sg13g2_decap_8
XFILLER_33_537 VPWR VGND sg13g2_decap_8
XFILLER_14_773 VPWR VGND sg13g2_decap_8
XFILLER_9_221 VPWR VGND sg13g2_decap_8
XFILLER_9_298 VPWR VGND sg13g2_decap_8
XFILLER_47_1008 VPWR VGND sg13g2_decap_8
XFILLER_37_832 VPWR VGND sg13g2_decap_8
XFILLER_24_515 VPWR VGND sg13g2_decap_8
XFILLER_34_19 VPWR VGND sg13g2_decap_8
XFILLER_36_375 VPWR VGND sg13g2_decap_8
XFILLER_20_754 VPWR VGND sg13g2_decap_8
XFILLER_28_876 VPWR VGND sg13g2_decap_8
XFILLER_43_824 VPWR VGND sg13g2_decap_8
XFILLER_15_504 VPWR VGND sg13g2_decap_8
XFILLER_27_364 VPWR VGND sg13g2_decap_8
XFILLER_42_334 VPWR VGND sg13g2_decap_8
XFILLER_11_732 VPWR VGND sg13g2_decap_8
XFILLER_23_592 VPWR VGND sg13g2_decap_8
XFILLER_24_74 VPWR VGND sg13g2_decap_8
XFILLER_10_242 VPWR VGND sg13g2_decap_8
XFILLER_7_714 VPWR VGND sg13g2_decap_8
XFILLER_6_235 VPWR VGND sg13g2_decap_8
X_094_ net31 _016_ _017_ VPWR VGND sg13g2_nand2_2
XFILLER_40_95 VPWR VGND sg13g2_decap_8
XFILLER_3_942 VPWR VGND sg13g2_decap_8
XFILLER_2_452 VPWR VGND sg13g2_decap_8
XFILLER_1_56 VPWR VGND sg13g2_decap_8
XFILLER_19_832 VPWR VGND sg13g2_decap_8
XFILLER_46_651 VPWR VGND sg13g2_decap_8
XFILLER_18_375 VPWR VGND sg13g2_decap_8
XFILLER_33_312 VPWR VGND sg13g2_decap_8
XFILLER_45_194 VPWR VGND sg13g2_decap_8
XFILLER_34_846 VPWR VGND sg13g2_decap_8
XFILLER_21_507 VPWR VGND sg13g2_decap_8
XFILLER_33_378 VPWR VGND sg13g2_decap_8
XFILLER_14_570 VPWR VGND sg13g2_decap_8
XFILLER_14_1018 VPWR VGND sg13g2_decap_8
XFILLER_46_0 VPWR VGND sg13g2_decap_8
XFILLER_25_824 VPWR VGND sg13g2_decap_8
XFILLER_24_334 VPWR VGND sg13g2_decap_4
XFILLER_36_194 VPWR VGND sg13g2_decap_8
XFILLER_12_529 VPWR VGND sg13g2_decap_8
XFILLER_40_838 VPWR VGND sg13g2_decap_8
XFILLER_20_551 VPWR VGND sg13g2_decap_8
XFILLER_4_739 VPWR VGND sg13g2_decap_8
XFILLER_10_32 VPWR VGND sg13g2_decap_8
XFILLER_3_249 VPWR VGND sg13g2_decap_8
XFILLER_0_945 VPWR VGND sg13g2_decap_8
XFILLER_48_938 VPWR VGND sg13g2_decap_8
XFILLER_19_74 VPWR VGND sg13g2_decap_8
XFILLER_47_448 VPWR VGND sg13g2_decap_8
XFILLER_27_161 VPWR VGND sg13g2_decap_8
XFILLER_28_673 VPWR VGND sg13g2_decap_8
XFILLER_43_621 VPWR VGND sg13g2_decap_8
XFILLER_16_846 VPWR VGND sg13g2_decap_8
XFILLER_35_40 VPWR VGND sg13g2_decap_8
XFILLER_37_1007 VPWR VGND sg13g2_decap_8
XFILLER_42_131 VPWR VGND sg13g2_decap_8
XFILLER_15_378 VPWR VGND sg13g2_decap_8
XFILLER_30_304 VPWR VGND sg13g2_decap_8
XFILLER_31_827 VPWR VGND sg13g2_decap_8
XFILLER_43_698 VPWR VGND sg13g2_decap_8
XFILLER_30_359 VPWR VGND sg13g2_decap_8
XFILLER_7_511 VPWR VGND sg13g2_decap_8
XFILLER_7_588 VPWR VGND sg13g2_decap_8
X_077_ mod1.i_out_8psk\[0\] _041_ net29 VPWR VGND sg13g2_and2_1
XFILLER_18_4 VPWR VGND sg13g2_decap_8
XFILLER_39_949 VPWR VGND sg13g2_decap_8
XFILLER_25_109 VPWR VGND sg13g2_decap_8
XFILLER_18_172 VPWR VGND sg13g2_decap_8
XFILLER_34_643 VPWR VGND sg13g2_decap_8
XFILLER_33_131 VPWR VGND sg13g2_decap_8
XFILLER_22_849 VPWR VGND sg13g2_decap_8
XFILLER_33_175 VPWR VGND sg13g2_decap_8
XFILLER_5_1005 VPWR VGND sg13g2_decap_8
XFILLER_45_908 VPWR VGND sg13g2_decap_8
XFILLER_29_459 VPWR VGND sg13g2_decap_8
XFILLER_38_960 VPWR VGND sg13g2_decap_8
XFILLER_44_418 VPWR VGND sg13g2_decap_8
XFILLER_16_109 VPWR VGND sg13g2_decap_8
XFILLER_25_621 VPWR VGND sg13g2_decap_8
XFILLER_13_816 VPWR VGND sg13g2_decap_8
XFILLER_9_809 VPWR VGND sg13g2_decap_8
XFILLER_12_326 VPWR VGND sg13g2_decap_8
XFILLER_24_186 VPWR VGND sg13g2_fill_2
XFILLER_25_698 VPWR VGND sg13g2_decap_8
XFILLER_40_635 VPWR VGND sg13g2_decap_8
XFILLER_8_319 VPWR VGND sg13g2_decap_8
XFILLER_21_871 VPWR VGND sg13g2_decap_8
XFILLER_21_53 VPWR VGND sg13g2_decap_8
XFILLER_4_536 VPWR VGND sg13g2_decap_8
XFILLER_0_742 VPWR VGND sg13g2_decap_8
XFILLER_48_735 VPWR VGND sg13g2_decap_8
XFILLER_47_245 VPWR VGND sg13g2_decap_8
XFILLER_16_643 VPWR VGND sg13g2_decap_8
XFILLER_28_470 VPWR VGND sg13g2_decap_8
XFILLER_44_985 VPWR VGND sg13g2_decap_8
XFILLER_43_495 VPWR VGND sg13g2_decap_8
XFILLER_31_624 VPWR VGND sg13g2_decap_8
XFILLER_30_145 VPWR VGND sg13g2_decap_8
XFILLER_12_893 VPWR VGND sg13g2_decap_8
XFILLER_8_886 VPWR VGND sg13g2_decap_8
XFILLER_7_77 VPWR VGND sg13g2_decap_8
XFILLER_7_385 VPWR VGND sg13g2_decap_8
X_129_ net14 VGND VPWR _007_ mod1.i_out_8psk\[1\] clknet_2_3__leaf_clk sg13g2_dfrbpq_1
XFILLER_39_746 VPWR VGND sg13g2_decap_8
XFILLER_38_256 VPWR VGND sg13g2_decap_8
XFILLER_35_941 VPWR VGND sg13g2_decap_8
XFILLER_34_440 VPWR VGND sg13g2_decap_8
XFILLER_42_19 VPWR VGND sg13g2_decap_8
XFILLER_21_123 VPWR VGND sg13g2_decap_8
XFILLER_22_646 VPWR VGND sg13g2_decap_8
XFILLER_1_539 VPWR VGND sg13g2_decap_8
XFILLER_45_705 VPWR VGND sg13g2_decap_8
XFILLER_29_278 VPWR VGND sg13g2_decap_8
XFILLER_44_215 VPWR VGND sg13g2_decap_8
XFILLER_29_289 VPWR VGND sg13g2_fill_2
XFILLER_16_53 VPWR VGND sg13g2_decap_8
XFILLER_26_952 VPWR VGND sg13g2_decap_8
XFILLER_41_922 VPWR VGND sg13g2_decap_8
XFILLER_13_613 VPWR VGND sg13g2_decap_8
XFILLER_25_495 VPWR VGND sg13g2_decap_8
XFILLER_9_606 VPWR VGND sg13g2_decap_8
XFILLER_12_123 VPWR VGND sg13g2_decap_8
XFILLER_40_432 VPWR VGND sg13g2_decap_8
XFILLER_41_999 VPWR VGND sg13g2_decap_8
XFILLER_8_116 VPWR VGND sg13g2_decap_8
XFILLER_5_823 VPWR VGND sg13g2_decap_8
XFILLER_32_96 VPWR VGND sg13g2_decap_8
XFILLER_4_333 VPWR VGND sg13g2_decap_8
XFILLER_48_532 VPWR VGND sg13g2_decap_8
XFILLER_16_440 VPWR VGND sg13g2_decap_8
XFILLER_17_952 VPWR VGND sg13g2_decap_8
XFILLER_35_248 VPWR VGND sg13g2_decap_8
XFILLER_44_782 VPWR VGND sg13g2_decap_8
XFILLER_32_922 VPWR VGND sg13g2_decap_8
XFILLER_43_292 VPWR VGND sg13g2_decap_8
XFILLER_31_421 VPWR VGND sg13g2_decap_8
XFILLER_32_999 VPWR VGND sg13g2_decap_8
XFILLER_12_690 VPWR VGND sg13g2_decap_8
XFILLER_31_498 VPWR VGND sg13g2_decap_8
XFILLER_8_683 VPWR VGND sg13g2_decap_8
XFILLER_7_182 VPWR VGND sg13g2_decap_8
XFILLER_39_543 VPWR VGND sg13g2_decap_8
XFILLER_2_1019 VPWR VGND sg13g2_decap_8
XFILLER_27_749 VPWR VGND sg13g2_decap_8
XFILLER_42_719 VPWR VGND sg13g2_decap_8
XFILLER_23_900 VPWR VGND sg13g2_decap_8
XFILLER_41_207 VPWR VGND sg13g2_decap_8
XFILLER_22_443 VPWR VGND sg13g2_decap_8
XFILLER_10_627 VPWR VGND sg13g2_decap_8
XFILLER_23_977 VPWR VGND sg13g2_decap_8
XFILLER_2_837 VPWR VGND sg13g2_decap_8
XFILLER_1_336 VPWR VGND sg13g2_decap_8
XFILLER_49_329 VPWR VGND sg13g2_decap_8
XFILLER_45_502 VPWR VGND sg13g2_decap_8
XFILLER_27_63 VPWR VGND sg13g2_decap_8
XFILLER_45_579 VPWR VGND sg13g2_decap_8
XFILLER_17_259 VPWR VGND sg13g2_decap_8
XFILLER_33_719 VPWR VGND sg13g2_decap_8
XFILLER_13_410 VPWR VGND sg13g2_decap_8
XFILLER_32_229 VPWR VGND sg13g2_decap_8
XFILLER_43_40 VPWR VGND sg13g2_decap_8
XFILLER_14_955 VPWR VGND sg13g2_decap_8
XFILLER_9_403 VPWR VGND sg13g2_decap_8
XFILLER_41_796 VPWR VGND sg13g2_decap_8
XFILLER_13_487 VPWR VGND sg13g2_decap_8
XFILLER_5_620 VPWR VGND sg13g2_decap_8
XFILLER_4_130 VPWR VGND sg13g2_decap_8
XFILLER_5_697 VPWR VGND sg13g2_decap_8
XFILLER_4_67 VPWR VGND sg13g2_decap_8
XFILLER_49_896 VPWR VGND sg13g2_decap_8
XFILLER_36_557 VPWR VGND sg13g2_decap_8
XFILLER_23_218 VPWR VGND sg13g2_decap_4
XFILLER_16_270 VPWR VGND sg13g2_decap_8
XFILLER_20_936 VPWR VGND sg13g2_decap_8
XFILLER_31_295 VPWR VGND sg13g2_decap_8
XFILLER_32_796 VPWR VGND sg13g2_decap_8
XFILLER_9_970 VPWR VGND sg13g2_decap_8
XFILLER_8_480 VPWR VGND sg13g2_decap_8
XFILLER_27_546 VPWR VGND sg13g2_decap_8
XFILLER_42_516 VPWR VGND sg13g2_decap_8
XFILLER_14_207 VPWR VGND sg13g2_decap_8
Xfanout11 _036_ net11 VPWR VGND sg13g2_buf_8
XFILLER_11_914 VPWR VGND sg13g2_decap_8
XFILLER_22_240 VPWR VGND sg13g2_decap_8
XFILLER_23_774 VPWR VGND sg13g2_decap_8
XFILLER_10_424 VPWR VGND sg13g2_decap_8
XFILLER_13_32 VPWR VGND sg13g2_decap_8
XFILLER_6_417 VPWR VGND sg13g2_decap_8
XFILLER_2_634 VPWR VGND sg13g2_decap_8
XFILLER_1_133 VPWR VGND sg13g2_decap_8
XFILLER_49_126 VPWR VGND sg13g2_decap_8
XFILLER_46_833 VPWR VGND sg13g2_decap_8
XFILLER_38_95 VPWR VGND sg13g2_decap_8
XFILLER_18_557 VPWR VGND sg13g2_decap_8
XFILLER_45_376 VPWR VGND sg13g2_decap_8
XFILLER_33_516 VPWR VGND sg13g2_decap_8
XFILLER_9_200 VPWR VGND sg13g2_decap_8
XFILLER_14_752 VPWR VGND sg13g2_decap_8
XFILLER_41_593 VPWR VGND sg13g2_decap_8
XFILLER_13_284 VPWR VGND sg13g2_decap_8
XFILLER_9_277 VPWR VGND sg13g2_decap_8
XFILLER_10_991 VPWR VGND sg13g2_decap_8
XFILLER_6_984 VPWR VGND sg13g2_decap_8
XFILLER_5_494 VPWR VGND sg13g2_decap_8
XFILLER_49_693 VPWR VGND sg13g2_decap_8
XFILLER_37_811 VPWR VGND sg13g2_decap_8
XFILLER_36_354 VPWR VGND sg13g2_decap_8
XFILLER_37_888 VPWR VGND sg13g2_decap_8
X_142__32 VPWR VGND net37 sg13g2_tiehi
XFILLER_20_733 VPWR VGND sg13g2_decap_8
XFILLER_32_593 VPWR VGND sg13g2_decap_8
XFILLER_30_1024 VPWR VGND sg13g2_decap_4
XFILLER_43_803 VPWR VGND sg13g2_decap_8
XFILLER_27_343 VPWR VGND sg13g2_decap_8
XFILLER_28_855 VPWR VGND sg13g2_decap_8
XFILLER_42_313 VPWR VGND sg13g2_decap_8
XFILLER_11_711 VPWR VGND sg13g2_decap_8
XFILLER_23_571 VPWR VGND sg13g2_decap_8
XFILLER_24_53 VPWR VGND sg13g2_decap_8
XFILLER_10_221 VPWR VGND sg13g2_decap_8
XFILLER_6_214 VPWR VGND sg13g2_decap_8
XFILLER_11_788 VPWR VGND sg13g2_decap_8
XFILLER_10_298 VPWR VGND sg13g2_decap_8
X_093_ _017_ mod1.q_out_qam16\[2\] net11 VPWR VGND sg13g2_nand2_1
XFILLER_3_921 VPWR VGND sg13g2_decap_8
XFILLER_40_74 VPWR VGND sg13g2_decap_8
XFILLER_2_431 VPWR VGND sg13g2_decap_8
XFILLER_3_998 VPWR VGND sg13g2_decap_8
XFILLER_1_35 VPWR VGND sg13g2_decap_8
XFILLER_19_811 VPWR VGND sg13g2_decap_8
XFILLER_46_630 VPWR VGND sg13g2_decap_8
XFILLER_18_354 VPWR VGND sg13g2_decap_8
XFILLER_19_888 VPWR VGND sg13g2_decap_8
XFILLER_34_825 VPWR VGND sg13g2_decap_8
XFILLER_45_173 VPWR VGND sg13g2_decap_8
XFILLER_42_880 VPWR VGND sg13g2_decap_8
XFILLER_41_390 VPWR VGND sg13g2_decap_8
XFILLER_6_781 VPWR VGND sg13g2_decap_8
XFILLER_5_291 VPWR VGND sg13g2_decap_8
Xinput1 ui_in[1] net1 VPWR VGND sg13g2_buf_2
XFILLER_49_490 VPWR VGND sg13g2_decap_8
XFILLER_45_19 VPWR VGND sg13g2_decap_8
XFILLER_25_803 VPWR VGND sg13g2_decap_8
XFILLER_37_685 VPWR VGND sg13g2_decap_8
XFILLER_24_313 VPWR VGND sg13g2_decap_8
XFILLER_36_173 VPWR VGND sg13g2_decap_8
XFILLER_12_508 VPWR VGND sg13g2_decap_8
XFILLER_40_817 VPWR VGND sg13g2_decap_8
XFILLER_33_880 VPWR VGND sg13g2_decap_8
XFILLER_20_530 VPWR VGND sg13g2_decap_8
XFILLER_32_390 VPWR VGND sg13g2_decap_8
XFILLER_10_11 VPWR VGND sg13g2_decap_8
XFILLER_4_718 VPWR VGND sg13g2_decap_8
XFILLER_3_228 VPWR VGND sg13g2_decap_8
XFILLER_10_88 VPWR VGND sg13g2_decap_8
XFILLER_0_924 VPWR VGND sg13g2_decap_8
XFILLER_48_917 VPWR VGND sg13g2_decap_8
XFILLER_47_427 VPWR VGND sg13g2_decap_8
XFILLER_19_53 VPWR VGND sg13g2_decap_8
XFILLER_28_652 VPWR VGND sg13g2_decap_8
XFILLER_43_600 VPWR VGND sg13g2_decap_8
XFILLER_15_302 VPWR VGND sg13g2_decap_8
XFILLER_16_825 VPWR VGND sg13g2_decap_8
XFILLER_27_140 VPWR VGND sg13g2_decap_8
XFILLER_42_110 VPWR VGND sg13g2_decap_8
XFILLER_43_677 VPWR VGND sg13g2_decap_8
XFILLER_15_357 VPWR VGND sg13g2_decap_8
XFILLER_31_806 VPWR VGND sg13g2_decap_8
XFILLER_42_187 VPWR VGND sg13g2_decap_8
XFILLER_35_96 VPWR VGND sg13g2_decap_8
XFILLER_11_585 VPWR VGND sg13g2_decap_8
XFILLER_7_567 VPWR VGND sg13g2_decap_8
X_076_ net5 net4 mod1.qam16_mod.i_level\[2\] VPWR VGND sg13g2_xor2_1
XFILLER_3_795 VPWR VGND sg13g2_decap_8
XFILLER_39_928 VPWR VGND sg13g2_decap_8
XFILLER_38_449 VPWR VGND sg13g2_decap_8
XFILLER_47_994 VPWR VGND sg13g2_decap_8
XFILLER_18_151 VPWR VGND sg13g2_decap_8
XFILLER_19_685 VPWR VGND sg13g2_decap_8
XFILLER_33_110 VPWR VGND sg13g2_decap_8
XFILLER_34_622 VPWR VGND sg13g2_decap_8
XFILLER_21_305 VPWR VGND sg13g2_decap_8
XFILLER_22_828 VPWR VGND sg13g2_decap_8
XFILLER_34_699 VPWR VGND sg13g2_decap_8
XFILLER_5_1028 VPWR VGND sg13g2_fill_1
XFILLER_29_438 VPWR VGND sg13g2_decap_8
XFILLER_25_600 VPWR VGND sg13g2_decap_8
XFILLER_37_482 VPWR VGND sg13g2_decap_8
XFILLER_25_677 VPWR VGND sg13g2_decap_8
XFILLER_12_305 VPWR VGND sg13g2_decap_8
XFILLER_24_165 VPWR VGND sg13g2_decap_8
XFILLER_40_614 VPWR VGND sg13g2_decap_8
XFILLER_21_850 VPWR VGND sg13g2_decap_8
XFILLER_4_515 VPWR VGND sg13g2_decap_8
XFILLER_21_32 VPWR VGND sg13g2_decap_8
XFILLER_0_721 VPWR VGND sg13g2_decap_8
XFILLER_48_714 VPWR VGND sg13g2_decap_8
XFILLER_0_798 VPWR VGND sg13g2_decap_8
XFILLER_47_224 VPWR VGND sg13g2_decap_8
XFILLER_46_84 VPWR VGND sg13g2_decap_8
XFILLER_16_622 VPWR VGND sg13g2_decap_8
XFILLER_44_964 VPWR VGND sg13g2_decap_8
XFILLER_43_474 VPWR VGND sg13g2_decap_8
XFILLER_15_165 VPWR VGND sg13g2_decap_8
XFILLER_15_176 VPWR VGND sg13g2_fill_2
XFILLER_16_699 VPWR VGND sg13g2_decap_8
XFILLER_31_603 VPWR VGND sg13g2_decap_8
XFILLER_30_124 VPWR VGND sg13g2_decap_8
XFILLER_12_872 VPWR VGND sg13g2_decap_8
XFILLER_8_865 VPWR VGND sg13g2_decap_8
XFILLER_11_382 VPWR VGND sg13g2_decap_8
XFILLER_7_364 VPWR VGND sg13g2_decap_8
XFILLER_7_56 VPWR VGND sg13g2_decap_8
X_128_ net13 VGND VPWR _006_ mod1.i_out_8psk\[0\] clknet_2_0__leaf_clk sg13g2_dfrbpq_1
X_059_ VPWR _034_ net6 VGND sg13g2_inv_1
XFILLER_3_592 VPWR VGND sg13g2_decap_8
XFILLER_39_725 VPWR VGND sg13g2_decap_8
XFILLER_38_235 VPWR VGND sg13g2_decap_8
XFILLER_47_791 VPWR VGND sg13g2_decap_8
XFILLER_19_482 VPWR VGND sg13g2_decap_8
XFILLER_35_920 VPWR VGND sg13g2_decap_8
XFILLER_21_102 VPWR VGND sg13g2_decap_8
XFILLER_22_625 VPWR VGND sg13g2_decap_8
XFILLER_35_997 VPWR VGND sg13g2_decap_8
XFILLER_10_809 VPWR VGND sg13g2_decap_8
XFILLER_34_496 VPWR VGND sg13g2_decap_8
XFILLER_1_518 VPWR VGND sg13g2_decap_8
XFILLER_29_257 VPWR VGND sg13g2_decap_8
XFILLER_26_931 VPWR VGND sg13g2_decap_8
XFILLER_41_901 VPWR VGND sg13g2_decap_8
XFILLER_16_32 VPWR VGND sg13g2_decap_8
XFILLER_12_102 VPWR VGND sg13g2_decap_8
XFILLER_25_474 VPWR VGND sg13g2_decap_8
XFILLER_40_411 VPWR VGND sg13g2_decap_8
XFILLER_41_978 VPWR VGND sg13g2_decap_8
XFILLER_13_669 VPWR VGND sg13g2_decap_8
XFILLER_12_179 VPWR VGND sg13g2_decap_8
XFILLER_40_488 VPWR VGND sg13g2_decap_8
XFILLER_5_802 VPWR VGND sg13g2_decap_8
XFILLER_32_75 VPWR VGND sg13g2_decap_8
XFILLER_4_312 VPWR VGND sg13g2_decap_8
XFILLER_5_879 VPWR VGND sg13g2_decap_8
XFILLER_4_389 VPWR VGND sg13g2_decap_8
XFILLER_48_511 VPWR VGND sg13g2_decap_8
XFILLER_0_595 VPWR VGND sg13g2_decap_8
XFILLER_48_588 VPWR VGND sg13g2_decap_8
XFILLER_17_931 VPWR VGND sg13g2_decap_8
XFILLER_36_739 VPWR VGND sg13g2_decap_8
XFILLER_28_290 VPWR VGND sg13g2_fill_2
XFILLER_32_901 VPWR VGND sg13g2_decap_8
XFILLER_44_761 VPWR VGND sg13g2_decap_8
XFILLER_31_400 VPWR VGND sg13g2_decap_8
XFILLER_43_271 VPWR VGND sg13g2_decap_8
XFILLER_16_496 VPWR VGND sg13g2_decap_8
XFILLER_31_477 VPWR VGND sg13g2_decap_8
XFILLER_32_978 VPWR VGND sg13g2_decap_8
XFILLER_8_662 VPWR VGND sg13g2_decap_8
XFILLER_7_161 VPWR VGND sg13g2_decap_8
XFILLER_39_522 VPWR VGND sg13g2_decap_8
XFILLER_27_728 VPWR VGND sg13g2_decap_8
XFILLER_39_599 VPWR VGND sg13g2_decap_8
XFILLER_19_290 VPWR VGND sg13g2_decap_8
XFILLER_22_422 VPWR VGND sg13g2_decap_8
XFILLER_23_956 VPWR VGND sg13g2_decap_8
XFILLER_35_794 VPWR VGND sg13g2_decap_8
XFILLER_10_606 VPWR VGND sg13g2_decap_8
XFILLER_22_499 VPWR VGND sg13g2_decap_8
XFILLER_5_109 VPWR VGND sg13g2_decap_8
XFILLER_2_816 VPWR VGND sg13g2_decap_8
XFILLER_1_315 VPWR VGND sg13g2_decap_8
XFILLER_49_308 VPWR VGND sg13g2_decap_8
XFILLER_18_739 VPWR VGND sg13g2_decap_8
XFILLER_27_42 VPWR VGND sg13g2_decap_8
XFILLER_45_558 VPWR VGND sg13g2_decap_8
XFILLER_17_238 VPWR VGND sg13g2_decap_8
XFILLER_32_208 VPWR VGND sg13g2_decap_8
XFILLER_14_934 VPWR VGND sg13g2_decap_8
XFILLER_41_775 VPWR VGND sg13g2_decap_8
XFILLER_13_466 VPWR VGND sg13g2_decap_8
XFILLER_43_96 VPWR VGND sg13g2_decap_8
XFILLER_9_459 VPWR VGND sg13g2_decap_8
XFILLER_5_676 VPWR VGND sg13g2_decap_8
XFILLER_4_186 VPWR VGND sg13g2_decap_8
XFILLER_4_46 VPWR VGND sg13g2_decap_8
XFILLER_1_882 VPWR VGND sg13g2_decap_8
XFILLER_49_875 VPWR VGND sg13g2_decap_8
XFILLER_0_392 VPWR VGND sg13g2_decap_8
XFILLER_48_385 VPWR VGND sg13g2_decap_8
XFILLER_36_536 VPWR VGND sg13g2_decap_8
XFILLER_20_915 VPWR VGND sg13g2_decap_8
XFILLER_32_775 VPWR VGND sg13g2_decap_8
XFILLER_31_274 VPWR VGND sg13g2_decap_8
XFILLER_27_525 VPWR VGND sg13g2_decap_8
XFILLER_39_396 VPWR VGND sg13g2_decap_8
Xfanout12 _036_ net12 VPWR VGND sg13g2_buf_1
XFILLER_35_591 VPWR VGND sg13g2_decap_8
XFILLER_23_753 VPWR VGND sg13g2_decap_8
XFILLER_10_403 VPWR VGND sg13g2_decap_8
XFILLER_13_11 VPWR VGND sg13g2_decap_8
XFILLER_13_88 VPWR VGND sg13g2_decap_8
XFILLER_2_613 VPWR VGND sg13g2_decap_8
XFILLER_8_4 VPWR VGND sg13g2_decap_8
XFILLER_1_112 VPWR VGND sg13g2_decap_8
XFILLER_49_105 VPWR VGND sg13g2_decap_8
XFILLER_1_189 VPWR VGND sg13g2_decap_8
XFILLER_46_812 VPWR VGND sg13g2_decap_8
XFILLER_38_74 VPWR VGND sg13g2_decap_8
XFILLER_18_536 VPWR VGND sg13g2_decap_8
XFILLER_46_889 VPWR VGND sg13g2_decap_8
XFILLER_45_355 VPWR VGND sg13g2_decap_8
XFILLER_14_731 VPWR VGND sg13g2_decap_8
XFILLER_41_572 VPWR VGND sg13g2_decap_8
XFILLER_13_263 VPWR VGND sg13g2_decap_8
XFILLER_9_256 VPWR VGND sg13g2_decap_8
XFILLER_10_970 VPWR VGND sg13g2_decap_8
XFILLER_6_963 VPWR VGND sg13g2_decap_8
XFILLER_5_473 VPWR VGND sg13g2_decap_8
XFILLER_49_672 VPWR VGND sg13g2_decap_8
XFILLER_48_182 VPWR VGND sg13g2_decap_8
XFILLER_36_333 VPWR VGND sg13g2_decap_8
XFILLER_37_867 VPWR VGND sg13g2_decap_8
XFILLER_20_712 VPWR VGND sg13g2_decap_8
XFILLER_32_572 VPWR VGND sg13g2_decap_8
XFILLER_20_789 VPWR VGND sg13g2_decap_8
XFILLER_30_1003 VPWR VGND sg13g2_decap_8
XFILLER_8_1026 VPWR VGND sg13g2_fill_2
XFILLER_47_609 VPWR VGND sg13g2_decap_8
XFILLER_46_119 VPWR VGND sg13g2_decap_8
XFILLER_28_834 VPWR VGND sg13g2_decap_8
XFILLER_27_322 VPWR VGND sg13g2_decap_8
XFILLER_39_193 VPWR VGND sg13g2_decap_8
XFILLER_43_859 VPWR VGND sg13g2_decap_8
XFILLER_15_539 VPWR VGND sg13g2_decap_8
XFILLER_27_399 VPWR VGND sg13g2_decap_8
XFILLER_42_369 VPWR VGND sg13g2_decap_8
XFILLER_23_550 VPWR VGND sg13g2_decap_8
XFILLER_24_32 VPWR VGND sg13g2_decap_8
XFILLER_10_200 VPWR VGND sg13g2_decap_8
XFILLER_11_767 VPWR VGND sg13g2_decap_8
XFILLER_10_277 VPWR VGND sg13g2_decap_8
XFILLER_7_749 VPWR VGND sg13g2_decap_8
X_092_ _016_ _045_ mod1.q_out_qpsk\[2\] _041_ mod1.psk8_mod.q_out\[2\] VPWR VGND sg13g2_a22oi_1
XFILLER_40_53 VPWR VGND sg13g2_decap_8
XFILLER_3_900 VPWR VGND sg13g2_decap_8
XFILLER_2_410 VPWR VGND sg13g2_decap_8
XFILLER_3_977 VPWR VGND sg13g2_decap_8
XFILLER_2_487 VPWR VGND sg13g2_decap_8
XFILLER_49_84 VPWR VGND sg13g2_decap_8
XFILLER_1_14 VPWR VGND sg13g2_decap_8
XFILLER_37_119 VPWR VGND sg13g2_decap_8
XFILLER_18_333 VPWR VGND sg13g2_decap_8
XFILLER_19_867 VPWR VGND sg13g2_decap_8
XFILLER_46_686 VPWR VGND sg13g2_decap_8
XFILLER_45_152 VPWR VGND sg13g2_decap_8
XFILLER_34_804 VPWR VGND sg13g2_decap_8
XFILLER_33_347 VPWR VGND sg13g2_decap_4
XFILLER_6_760 VPWR VGND sg13g2_decap_8
XFILLER_5_270 VPWR VGND sg13g2_decap_8
Xinput2 ui_in[2] net2 VPWR VGND sg13g2_buf_2
XFILLER_36_152 VPWR VGND sg13g2_decap_8
XFILLER_37_664 VPWR VGND sg13g2_decap_8
XFILLER_25_859 VPWR VGND sg13g2_decap_8
XFILLER_24_358 VPWR VGND sg13g2_decap_8
XFILLER_20_586 VPWR VGND sg13g2_decap_8
XFILLER_3_207 VPWR VGND sg13g2_decap_8
XFILLER_10_67 VPWR VGND sg13g2_decap_8
XFILLER_0_903 VPWR VGND sg13g2_decap_8
XFILLER_47_406 VPWR VGND sg13g2_decap_8
XFILLER_19_32 VPWR VGND sg13g2_decap_8
XFILLER_28_631 VPWR VGND sg13g2_decap_8
XFILLER_16_804 VPWR VGND sg13g2_decap_8
XFILLER_43_656 VPWR VGND sg13g2_decap_8
XFILLER_27_196 VPWR VGND sg13g2_decap_8
XFILLER_35_75 VPWR VGND sg13g2_decap_8
XFILLER_42_166 VPWR VGND sg13g2_decap_8
XFILLER_11_564 VPWR VGND sg13g2_decap_8
XFILLER_7_546 VPWR VGND sg13g2_decap_8
X_075_ Demo1.qam16_bits\[3\] net11 net24 VPWR VGND sg13g2_and2_1
XFILLER_3_774 VPWR VGND sg13g2_decap_8
XFILLER_2_284 VPWR VGND sg13g2_decap_8
XFILLER_39_907 VPWR VGND sg13g2_decap_8
XFILLER_38_428 VPWR VGND sg13g2_decap_8
XFILLER_20_1013 VPWR VGND sg13g2_decap_8
XFILLER_47_973 VPWR VGND sg13g2_decap_8
XFILLER_18_130 VPWR VGND sg13g2_decap_8
XFILLER_19_664 VPWR VGND sg13g2_decap_8
XFILLER_34_601 VPWR VGND sg13g2_decap_8
XFILLER_46_483 VPWR VGND sg13g2_decap_8
XFILLER_22_807 VPWR VGND sg13g2_decap_8
XFILLER_34_678 VPWR VGND sg13g2_decap_8
XFILLER_30_884 VPWR VGND sg13g2_decap_8
XFILLER_29_417 VPWR VGND sg13g2_decap_8
XFILLER_37_461 VPWR VGND sg13g2_decap_8
XFILLER_38_995 VPWR VGND sg13g2_decap_8
XFILLER_24_144 VPWR VGND sg13g2_decap_8
XFILLER_25_656 VPWR VGND sg13g2_decap_8
XFILLER_24_188 VPWR VGND sg13g2_fill_1
XFILLER_20_372 VPWR VGND sg13g2_decap_8
XFILLER_21_11 VPWR VGND sg13g2_decap_8
XFILLER_21_88 VPWR VGND sg13g2_decap_8
XFILLER_0_700 VPWR VGND sg13g2_decap_8
XFILLER_43_1013 VPWR VGND sg13g2_decap_8
XFILLER_47_203 VPWR VGND sg13g2_decap_8
XFILLER_0_777 VPWR VGND sg13g2_decap_8
XFILLER_29_984 VPWR VGND sg13g2_decap_8
XFILLER_35_409 VPWR VGND sg13g2_decap_8
XFILLER_46_63 VPWR VGND sg13g2_decap_8
XFILLER_44_943 VPWR VGND sg13g2_decap_8
XFILLER_16_601 VPWR VGND sg13g2_decap_8
XFILLER_43_453 VPWR VGND sg13g2_decap_8
XFILLER_15_144 VPWR VGND sg13g2_decap_8
XFILLER_16_678 VPWR VGND sg13g2_decap_8
XFILLER_30_103 VPWR VGND sg13g2_decap_8
XFILLER_31_659 VPWR VGND sg13g2_decap_8
XFILLER_12_851 VPWR VGND sg13g2_decap_8
XFILLER_8_844 VPWR VGND sg13g2_decap_8
XFILLER_7_35 VPWR VGND sg13g2_decap_8
XFILLER_11_361 VPWR VGND sg13g2_decap_8
XFILLER_7_343 VPWR VGND sg13g2_decap_8
X_127_ net13 VGND VPWR _010_ mod1.psk8_mod.q_out\[2\] clknet_2_0__leaf_clk sg13g2_dfrbpq_1
X_058_ VPWR _033_ net7 VGND sg13g2_inv_1
XFILLER_3_571 VPWR VGND sg13g2_decap_8
XFILLER_30_5 VPWR VGND sg13g2_decap_8
XFILLER_23_4 VPWR VGND sg13g2_decap_8
XFILLER_39_704 VPWR VGND sg13g2_decap_8
XFILLER_38_214 VPWR VGND sg13g2_decap_8
XFILLER_47_770 VPWR VGND sg13g2_decap_8
XFILLER_19_461 VPWR VGND sg13g2_decap_8
XFILLER_46_280 VPWR VGND sg13g2_decap_8
XFILLER_35_976 VPWR VGND sg13g2_decap_8
XFILLER_22_604 VPWR VGND sg13g2_decap_8
XFILLER_34_475 VPWR VGND sg13g2_decap_8
XFILLER_21_169 VPWR VGND sg13g2_decap_8
XFILLER_30_681 VPWR VGND sg13g2_decap_8
XFILLER_27_1008 VPWR VGND sg13g2_decap_8
XFILLER_29_236 VPWR VGND sg13g2_decap_8
XFILLER_16_11 VPWR VGND sg13g2_decap_8
XFILLER_26_910 VPWR VGND sg13g2_decap_8
XFILLER_38_792 VPWR VGND sg13g2_decap_8
XFILLER_25_453 VPWR VGND sg13g2_decap_8
XFILLER_26_987 VPWR VGND sg13g2_decap_8
XFILLER_41_957 VPWR VGND sg13g2_decap_8
XFILLER_13_648 VPWR VGND sg13g2_decap_8
XFILLER_16_88 VPWR VGND sg13g2_decap_8
XFILLER_12_158 VPWR VGND sg13g2_decap_8
XFILLER_40_467 VPWR VGND sg13g2_decap_8
XFILLER_32_54 VPWR VGND sg13g2_decap_8
XFILLER_10_1012 VPWR VGND sg13g2_decap_8
XFILLER_5_858 VPWR VGND sg13g2_decap_8
XFILLER_4_368 VPWR VGND sg13g2_decap_8
XFILLER_0_574 VPWR VGND sg13g2_decap_8
XFILLER_48_567 VPWR VGND sg13g2_decap_8
XFILLER_36_718 VPWR VGND sg13g2_decap_8
XFILLER_17_910 VPWR VGND sg13g2_decap_8
XFILLER_29_781 VPWR VGND sg13g2_decap_8
XFILLER_35_228 VPWR VGND sg13g2_decap_8
XFILLER_44_740 VPWR VGND sg13g2_decap_8
XFILLER_43_250 VPWR VGND sg13g2_decap_8
XFILLER_16_475 VPWR VGND sg13g2_decap_8
XFILLER_17_987 VPWR VGND sg13g2_decap_8
XFILLER_32_957 VPWR VGND sg13g2_decap_8
XFILLER_31_456 VPWR VGND sg13g2_decap_8
XFILLER_8_641 VPWR VGND sg13g2_decap_8
XFILLER_7_140 VPWR VGND sg13g2_decap_8
XFILLER_39_501 VPWR VGND sg13g2_decap_8
XFILLER_27_707 VPWR VGND sg13g2_decap_8
XFILLER_39_578 VPWR VGND sg13g2_decap_8
XFILLER_26_228 VPWR VGND sg13g2_fill_1
XFILLER_26_239 VPWR VGND sg13g2_decap_8
XFILLER_22_401 VPWR VGND sg13g2_decap_8
XFILLER_35_773 VPWR VGND sg13g2_decap_8
XFILLER_23_935 VPWR VGND sg13g2_decap_8
XFILLER_34_294 VPWR VGND sg13g2_decap_4
XFILLER_22_478 VPWR VGND sg13g2_decap_8
XFILLER_18_718 VPWR VGND sg13g2_decap_8
XFILLER_40_1027 VPWR VGND sg13g2_fill_2
XFILLER_45_537 VPWR VGND sg13g2_decap_8
XFILLER_17_217 VPWR VGND sg13g2_decap_8
XFILLER_27_21 VPWR VGND sg13g2_decap_8
XFILLER_14_913 VPWR VGND sg13g2_decap_8
XFILLER_26_784 VPWR VGND sg13g2_decap_8
XFILLER_27_98 VPWR VGND sg13g2_decap_8
XFILLER_25_283 VPWR VGND sg13g2_decap_8
XFILLER_41_754 VPWR VGND sg13g2_decap_8
XFILLER_13_445 VPWR VGND sg13g2_decap_8
XFILLER_43_75 VPWR VGND sg13g2_decap_8
XFILLER_9_438 VPWR VGND sg13g2_decap_8
XFILLER_40_264 VPWR VGND sg13g2_decap_8
XFILLER_5_655 VPWR VGND sg13g2_decap_8
XFILLER_4_165 VPWR VGND sg13g2_decap_8
XFILLER_4_25 VPWR VGND sg13g2_decap_8
XFILLER_1_861 VPWR VGND sg13g2_decap_8
XFILLER_0_371 VPWR VGND sg13g2_decap_8
XFILLER_49_854 VPWR VGND sg13g2_decap_8
XFILLER_48_364 VPWR VGND sg13g2_decap_8
XFILLER_36_515 VPWR VGND sg13g2_decap_8
XFILLER_17_784 VPWR VGND sg13g2_decap_8
XFILLER_31_253 VPWR VGND sg13g2_decap_8
XFILLER_32_754 VPWR VGND sg13g2_decap_8
XFILLER_27_504 VPWR VGND sg13g2_decap_8
XFILLER_39_375 VPWR VGND sg13g2_decap_8
Xfanout13 net15 net13 VPWR VGND sg13g2_buf_8
XFILLER_23_732 VPWR VGND sg13g2_decap_8
XFILLER_35_570 VPWR VGND sg13g2_decap_8
XFILLER_11_949 VPWR VGND sg13g2_decap_8
XFILLER_10_459 VPWR VGND sg13g2_decap_8
XFILLER_13_67 VPWR VGND sg13g2_decap_8
XFILLER_2_669 VPWR VGND sg13g2_decap_8
XFILLER_1_168 VPWR VGND sg13g2_decap_8
XFILLER_38_53 VPWR VGND sg13g2_decap_8
XFILLER_18_515 VPWR VGND sg13g2_decap_8
XFILLER_46_868 VPWR VGND sg13g2_decap_8
XFILLER_45_334 VPWR VGND sg13g2_decap_8
XFILLER_14_710 VPWR VGND sg13g2_decap_8
XFILLER_26_581 VPWR VGND sg13g2_decap_8
XFILLER_41_551 VPWR VGND sg13g2_decap_8
XFILLER_13_242 VPWR VGND sg13g2_decap_8
XFILLER_14_787 VPWR VGND sg13g2_decap_8
XFILLER_9_235 VPWR VGND sg13g2_decap_8
XFILLER_6_942 VPWR VGND sg13g2_decap_8
XFILLER_5_452 VPWR VGND sg13g2_decap_8
XFILLER_49_651 VPWR VGND sg13g2_decap_8
XFILLER_48_161 VPWR VGND sg13g2_decap_8
XFILLER_36_312 VPWR VGND sg13g2_decap_8
XFILLER_37_846 VPWR VGND sg13g2_decap_8
XFILLER_17_581 VPWR VGND sg13g2_decap_8
XFILLER_24_529 VPWR VGND sg13g2_decap_8
XFILLER_36_389 VPWR VGND sg13g2_decap_8
XFILLER_32_551 VPWR VGND sg13g2_decap_8
XFILLER_20_768 VPWR VGND sg13g2_decap_8
XFILLER_8_1005 VPWR VGND sg13g2_decap_8
XFILLER_27_301 VPWR VGND sg13g2_decap_8
XFILLER_28_813 VPWR VGND sg13g2_decap_8
XFILLER_39_172 VPWR VGND sg13g2_decap_8
XFILLER_15_518 VPWR VGND sg13g2_decap_8
XFILLER_27_378 VPWR VGND sg13g2_decap_8
XFILLER_43_838 VPWR VGND sg13g2_decap_8
XFILLER_42_348 VPWR VGND sg13g2_decap_8
XFILLER_24_11 VPWR VGND sg13g2_decap_8
XFILLER_11_746 VPWR VGND sg13g2_decap_8
XFILLER_24_88 VPWR VGND sg13g2_decap_8
XFILLER_10_256 VPWR VGND sg13g2_decap_8
XFILLER_7_728 VPWR VGND sg13g2_decap_8
XFILLER_6_249 VPWR VGND sg13g2_decap_8
X_091_ net30 _046_ _015_ VPWR VGND sg13g2_nand2_2
XFILLER_40_32 VPWR VGND sg13g2_decap_8
XFILLER_3_956 VPWR VGND sg13g2_decap_8
XFILLER_46_1022 VPWR VGND sg13g2_decap_8
XFILLER_2_466 VPWR VGND sg13g2_decap_8
XFILLER_49_63 VPWR VGND sg13g2_decap_8
XFILLER_18_312 VPWR VGND sg13g2_decap_8
XFILLER_19_846 VPWR VGND sg13g2_decap_8
XFILLER_46_665 VPWR VGND sg13g2_decap_8
XFILLER_45_131 VPWR VGND sg13g2_decap_8
XFILLER_18_389 VPWR VGND sg13g2_decap_8
XFILLER_33_326 VPWR VGND sg13g2_decap_8
XFILLER_14_584 VPWR VGND sg13g2_decap_8
XFILLER_28_109 VPWR VGND sg13g2_decap_8
Xinput3 ui_in[3] net3 VPWR VGND sg13g2_buf_2
XFILLER_37_643 VPWR VGND sg13g2_decap_8
XFILLER_36_131 VPWR VGND sg13g2_decap_8
XFILLER_25_838 VPWR VGND sg13g2_decap_8
XFILLER_20_565 VPWR VGND sg13g2_decap_8
XFILLER_10_46 VPWR VGND sg13g2_decap_8
XFILLER_0_959 VPWR VGND sg13g2_decap_8
XFILLER_19_11 VPWR VGND sg13g2_decap_8
XFILLER_19_109 VPWR VGND sg13g2_decap_8
XFILLER_19_88 VPWR VGND sg13g2_decap_8
XFILLER_28_610 VPWR VGND sg13g2_decap_8
XFILLER_43_635 VPWR VGND sg13g2_decap_8
XFILLER_27_175 VPWR VGND sg13g2_decap_8
XFILLER_28_687 VPWR VGND sg13g2_decap_8
XFILLER_42_145 VPWR VGND sg13g2_decap_8
XFILLER_35_54 VPWR VGND sg13g2_decap_8
XFILLER_30_318 VPWR VGND sg13g2_decap_8
XFILLER_24_893 VPWR VGND sg13g2_decap_8
XFILLER_11_543 VPWR VGND sg13g2_decap_8
XFILLER_7_525 VPWR VGND sg13g2_decap_8
X_143_ net14 VGND VPWR _000_ mod1.bpsk_mod.i_out\[2\] clknet_2_0__leaf_clk sg13g2_dfrbpq_1
X_074_ net23 _044_ VPWR VGND sg13g2_inv_2
XFILLER_3_753 VPWR VGND sg13g2_decap_8
XFILLER_2_263 VPWR VGND sg13g2_decap_8
XFILLER_38_407 VPWR VGND sg13g2_decap_8
XFILLER_47_952 VPWR VGND sg13g2_decap_8
XFILLER_19_643 VPWR VGND sg13g2_decap_8
XFILLER_46_462 VPWR VGND sg13g2_decap_8
XFILLER_18_186 VPWR VGND sg13g2_decap_8
XFILLER_33_145 VPWR VGND sg13g2_fill_2
XFILLER_34_657 VPWR VGND sg13g2_decap_8
XFILLER_15_882 VPWR VGND sg13g2_decap_8
XFILLER_14_381 VPWR VGND sg13g2_decap_8
XFILLER_33_189 VPWR VGND sg13g2_decap_8
XFILLER_30_863 VPWR VGND sg13g2_decap_8
XFILLER_5_1019 VPWR VGND sg13g2_decap_8
XFILLER_37_440 VPWR VGND sg13g2_decap_8
XFILLER_38_974 VPWR VGND sg13g2_decap_8
XFILLER_24_123 VPWR VGND sg13g2_decap_8
XFILLER_25_635 VPWR VGND sg13g2_decap_8
XFILLER_40_649 VPWR VGND sg13g2_decap_8
XFILLER_20_340 VPWR VGND sg13g2_decap_4
XFILLER_20_351 VPWR VGND sg13g2_decap_8
XFILLER_20_384 VPWR VGND sg13g2_decap_8
XFILLER_21_885 VPWR VGND sg13g2_decap_8
XFILLER_21_67 VPWR VGND sg13g2_decap_8
XFILLER_0_756 VPWR VGND sg13g2_decap_8
XFILLER_48_749 VPWR VGND sg13g2_decap_8
XFILLER_47_259 VPWR VGND sg13g2_decap_8
XFILLER_46_42 VPWR VGND sg13g2_decap_8
XFILLER_29_963 VPWR VGND sg13g2_decap_8
XFILLER_44_922 VPWR VGND sg13g2_decap_8
XFILLER_28_484 VPWR VGND sg13g2_decap_8
XFILLER_43_432 VPWR VGND sg13g2_decap_8
XFILLER_15_123 VPWR VGND sg13g2_decap_8
XFILLER_16_657 VPWR VGND sg13g2_decap_8
XFILLER_44_999 VPWR VGND sg13g2_decap_8
XFILLER_12_830 VPWR VGND sg13g2_decap_8
XFILLER_24_690 VPWR VGND sg13g2_decap_8
XFILLER_31_638 VPWR VGND sg13g2_decap_8
XFILLER_8_823 VPWR VGND sg13g2_decap_8
XFILLER_11_340 VPWR VGND sg13g2_decap_8
XFILLER_30_159 VPWR VGND sg13g2_decap_8
XFILLER_7_322 VPWR VGND sg13g2_decap_8
XFILLER_7_14 VPWR VGND sg13g2_decap_8
X_126_ net13 VGND VPWR _009_ mod1.psk8_mod.q_out\[1\] clknet_2_2__leaf_clk sg13g2_dfrbpq_1
XFILLER_7_399 VPWR VGND sg13g2_decap_8
X_057_ net5 mod1.qam16_mod.i_level\[3\] VPWR VGND sg13g2_inv_4
XFILLER_3_550 VPWR VGND sg13g2_decap_8
XFILLER_16_4 VPWR VGND sg13g2_decap_8
XFILLER_19_440 VPWR VGND sg13g2_decap_8
XFILLER_35_955 VPWR VGND sg13g2_decap_8
XFILLER_34_454 VPWR VGND sg13g2_decap_8
XFILLER_21_137 VPWR VGND sg13g2_decap_8
XFILLER_30_660 VPWR VGND sg13g2_decap_8
XFILLER_45_719 VPWR VGND sg13g2_decap_8
XFILLER_44_229 VPWR VGND sg13g2_decap_8
XFILLER_38_771 VPWR VGND sg13g2_decap_8
XFILLER_25_432 VPWR VGND sg13g2_decap_8
XFILLER_26_966 VPWR VGND sg13g2_decap_8
XFILLER_37_292 VPWR VGND sg13g2_decap_8
XFILLER_16_67 VPWR VGND sg13g2_decap_8
XFILLER_41_936 VPWR VGND sg13g2_decap_8
XFILLER_13_627 VPWR VGND sg13g2_decap_8
XFILLER_12_137 VPWR VGND sg13g2_decap_8
XFILLER_40_446 VPWR VGND sg13g2_decap_8
XFILLER_21_682 VPWR VGND sg13g2_decap_8
XFILLER_32_33 VPWR VGND sg13g2_decap_8
XFILLER_5_837 VPWR VGND sg13g2_decap_8
XFILLER_4_347 VPWR VGND sg13g2_decap_8
XFILLER_0_553 VPWR VGND sg13g2_decap_8
XFILLER_48_546 VPWR VGND sg13g2_decap_8
XFILLER_29_760 VPWR VGND sg13g2_decap_8
XFILLER_35_207 VPWR VGND sg13g2_decap_8
XFILLER_17_966 VPWR VGND sg13g2_decap_8
XFILLER_16_454 VPWR VGND sg13g2_decap_8
XFILLER_44_796 VPWR VGND sg13g2_decap_8
XFILLER_31_435 VPWR VGND sg13g2_decap_8
XFILLER_32_936 VPWR VGND sg13g2_decap_8
XFILLER_8_620 VPWR VGND sg13g2_decap_8
XFILLER_8_697 VPWR VGND sg13g2_decap_8
XFILLER_7_196 VPWR VGND sg13g2_decap_8
X_109_ VGND VPWR _024_ net1 net17 sg13g2_or2_1
XFILLER_39_557 VPWR VGND sg13g2_decap_8
XFILLER_26_207 VPWR VGND sg13g2_decap_8
XFILLER_23_914 VPWR VGND sg13g2_decap_8
XFILLER_35_752 VPWR VGND sg13g2_decap_8
XFILLER_34_273 VPWR VGND sg13g2_decap_8
XFILLER_22_457 VPWR VGND sg13g2_decap_8
XFILLER_33_1013 VPWR VGND sg13g2_decap_8
XFILLER_40_1006 VPWR VGND sg13g2_decap_8
XFILLER_45_516 VPWR VGND sg13g2_decap_8
XFILLER_27_77 VPWR VGND sg13g2_decap_8
XFILLER_26_763 VPWR VGND sg13g2_decap_8
XFILLER_41_733 VPWR VGND sg13g2_decap_8
XFILLER_13_424 VPWR VGND sg13g2_decap_8
XFILLER_25_262 VPWR VGND sg13g2_decap_8
XFILLER_43_54 VPWR VGND sg13g2_decap_8
XFILLER_9_417 VPWR VGND sg13g2_decap_8
XFILLER_14_969 VPWR VGND sg13g2_decap_8
XFILLER_40_243 VPWR VGND sg13g2_decap_8
XFILLER_5_634 VPWR VGND sg13g2_decap_8
XFILLER_4_144 VPWR VGND sg13g2_decap_8
XFILLER_1_840 VPWR VGND sg13g2_decap_8
XFILLER_49_833 VPWR VGND sg13g2_decap_8
XFILLER_0_350 VPWR VGND sg13g2_decap_8
XFILLER_48_343 VPWR VGND sg13g2_decap_8
XFILLER_1_1022 VPWR VGND sg13g2_decap_8
XFILLER_17_763 VPWR VGND sg13g2_decap_8
XFILLER_44_593 VPWR VGND sg13g2_decap_8
XFILLER_16_284 VPWR VGND sg13g2_decap_8
XFILLER_32_733 VPWR VGND sg13g2_decap_8
XFILLER_17_1008 VPWR VGND sg13g2_decap_8
XFILLER_13_991 VPWR VGND sg13g2_decap_8
XFILLER_9_984 VPWR VGND sg13g2_decap_8
XFILLER_8_494 VPWR VGND sg13g2_decap_8
XFILLER_39_332 VPWR VGND sg13g2_fill_2
XFILLER_23_711 VPWR VGND sg13g2_decap_8
Xfanout14 net15 net14 VPWR VGND sg13g2_buf_8
XFILLER_11_928 VPWR VGND sg13g2_decap_8
XFILLER_22_254 VPWR VGND sg13g2_decap_8
XFILLER_23_788 VPWR VGND sg13g2_decap_8
XFILLER_10_438 VPWR VGND sg13g2_decap_8
XFILLER_13_46 VPWR VGND sg13g2_decap_8
XFILLER_2_648 VPWR VGND sg13g2_decap_8
XFILLER_1_147 VPWR VGND sg13g2_decap_8
XFILLER_38_32 VPWR VGND sg13g2_decap_8
XFILLER_46_847 VPWR VGND sg13g2_decap_8
XFILLER_45_313 VPWR VGND sg13g2_decap_8
XFILLER_26_560 VPWR VGND sg13g2_decap_8
XFILLER_41_530 VPWR VGND sg13g2_decap_8
XFILLER_13_221 VPWR VGND sg13g2_decap_8
XFILLER_14_766 VPWR VGND sg13g2_decap_8
XFILLER_9_214 VPWR VGND sg13g2_decap_8
XFILLER_13_298 VPWR VGND sg13g2_decap_8
XFILLER_6_921 VPWR VGND sg13g2_decap_8
XFILLER_5_431 VPWR VGND sg13g2_decap_8
XFILLER_6_998 VPWR VGND sg13g2_decap_8
XFILLER_48_7 VPWR VGND sg13g2_decap_8
XFILLER_49_630 VPWR VGND sg13g2_decap_8
XFILLER_23_1012 VPWR VGND sg13g2_decap_8
XFILLER_48_140 VPWR VGND sg13g2_decap_8
XFILLER_37_825 VPWR VGND sg13g2_decap_8
XFILLER_24_508 VPWR VGND sg13g2_decap_8
XFILLER_36_368 VPWR VGND sg13g2_decap_8
XFILLER_45_880 VPWR VGND sg13g2_decap_8
XFILLER_17_560 VPWR VGND sg13g2_decap_8
XFILLER_44_390 VPWR VGND sg13g2_decap_8
XFILLER_32_530 VPWR VGND sg13g2_decap_8
XFILLER_20_747 VPWR VGND sg13g2_decap_8
XFILLER_9_781 VPWR VGND sg13g2_decap_8
XFILLER_8_291 VPWR VGND sg13g2_decap_8
XFILLER_8_1028 VPWR VGND sg13g2_fill_1
XFILLER_39_151 VPWR VGND sg13g2_decap_8
XFILLER_43_817 VPWR VGND sg13g2_decap_8
XFILLER_27_357 VPWR VGND sg13g2_decap_8
XFILLER_28_869 VPWR VGND sg13g2_decap_8
XFILLER_42_327 VPWR VGND sg13g2_decap_8
XFILLER_11_725 VPWR VGND sg13g2_decap_8
XFILLER_24_67 VPWR VGND sg13g2_decap_8
XFILLER_7_707 VPWR VGND sg13g2_decap_8
XFILLER_23_585 VPWR VGND sg13g2_decap_8
XFILLER_10_235 VPWR VGND sg13g2_decap_8
X_090_ _015_ mod1.psk8_mod.q_out\[1\] _041_ VPWR VGND sg13g2_nand2_1
XFILLER_40_11 VPWR VGND sg13g2_decap_8
XFILLER_6_228 VPWR VGND sg13g2_decap_8
XFILLER_3_935 VPWR VGND sg13g2_decap_8
XFILLER_40_88 VPWR VGND sg13g2_decap_8
XFILLER_46_1001 VPWR VGND sg13g2_decap_8
XFILLER_2_445 VPWR VGND sg13g2_decap_8
XFILLER_49_42 VPWR VGND sg13g2_decap_8
XFILLER_19_825 VPWR VGND sg13g2_decap_8
XFILLER_46_644 VPWR VGND sg13g2_decap_8
XFILLER_45_110 VPWR VGND sg13g2_decap_8
XFILLER_1_49 VPWR VGND sg13g2_decap_8
XFILLER_18_368 VPWR VGND sg13g2_decap_8
XFILLER_45_187 VPWR VGND sg13g2_decap_8
XFILLER_33_305 VPWR VGND sg13g2_decap_8
XFILLER_34_839 VPWR VGND sg13g2_decap_8
XFILLER_14_563 VPWR VGND sg13g2_decap_8
XFILLER_42_894 VPWR VGND sg13g2_decap_8
XFILLER_6_795 VPWR VGND sg13g2_decap_8
Xinput4 ui_in[4] net4 VPWR VGND sg13g2_buf_2
XFILLER_36_110 VPWR VGND sg13g2_decap_8
XFILLER_37_622 VPWR VGND sg13g2_decap_8
XFILLER_25_817 VPWR VGND sg13g2_decap_8
XFILLER_24_327 VPWR VGND sg13g2_decap_8
Xclkbuf_2_1__f_clk clknet_0_clk clknet_2_1__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_36_187 VPWR VGND sg13g2_decap_8
XFILLER_37_699 VPWR VGND sg13g2_decap_8
XFILLER_33_894 VPWR VGND sg13g2_decap_8
XFILLER_20_544 VPWR VGND sg13g2_decap_8
XFILLER_10_25 VPWR VGND sg13g2_decap_8
XFILLER_0_938 VPWR VGND sg13g2_decap_8
XFILLER_19_67 VPWR VGND sg13g2_decap_8
XFILLER_28_666 VPWR VGND sg13g2_decap_8
XFILLER_43_614 VPWR VGND sg13g2_decap_8
XFILLER_16_839 VPWR VGND sg13g2_decap_8
XFILLER_27_154 VPWR VGND sg13g2_decap_8
XFILLER_35_33 VPWR VGND sg13g2_decap_8
XFILLER_42_124 VPWR VGND sg13g2_decap_8
XFILLER_24_872 VPWR VGND sg13g2_decap_8
XFILLER_11_522 VPWR VGND sg13g2_decap_8
XFILLER_23_382 VPWR VGND sg13g2_decap_8
XFILLER_7_504 VPWR VGND sg13g2_decap_8
X_142_ net13 VGND VPWR net37 Demo1.qam16_bits\[3\] clknet_2_2__leaf_clk sg13g2_dfrbpq_2
XFILLER_11_599 VPWR VGND sg13g2_decap_8
X_073_ _044_ _041_ Demo1.epsk_de1.bit_out\[2\] net12 Demo1.qam16_bits\[2\] VPWR VGND
+ sg13g2_a22oi_1
XFILLER_3_732 VPWR VGND sg13g2_decap_8
XFILLER_2_242 VPWR VGND sg13g2_decap_8
XFILLER_47_931 VPWR VGND sg13g2_decap_8
XFILLER_19_622 VPWR VGND sg13g2_decap_8
XFILLER_46_441 VPWR VGND sg13g2_decap_8
XFILLER_18_165 VPWR VGND sg13g2_decap_8
XFILLER_19_699 VPWR VGND sg13g2_decap_8
XFILLER_33_124 VPWR VGND sg13g2_decap_8
XFILLER_34_636 VPWR VGND sg13g2_decap_8
XFILLER_15_861 VPWR VGND sg13g2_decap_8
XFILLER_21_319 VPWR VGND sg13g2_fill_1
XFILLER_42_691 VPWR VGND sg13g2_decap_8
XFILLER_14_360 VPWR VGND sg13g2_decap_8
XFILLER_30_842 VPWR VGND sg13g2_decap_8
XFILLER_6_592 VPWR VGND sg13g2_decap_8
XFILLER_37_0 VPWR VGND sg13g2_decap_8
XFILLER_2_81 VPWR VGND sg13g2_decap_8
XFILLER_38_953 VPWR VGND sg13g2_decap_8
XFILLER_24_102 VPWR VGND sg13g2_decap_8
XFILLER_25_614 VPWR VGND sg13g2_decap_8
XFILLER_37_496 VPWR VGND sg13g2_decap_8
XFILLER_13_809 VPWR VGND sg13g2_decap_8
XFILLER_12_319 VPWR VGND sg13g2_decap_8
XFILLER_24_179 VPWR VGND sg13g2_decap_8
XFILLER_33_691 VPWR VGND sg13g2_decap_8
XFILLER_40_628 VPWR VGND sg13g2_decap_8
XFILLER_21_864 VPWR VGND sg13g2_decap_8
XFILLER_21_46 VPWR VGND sg13g2_decap_8
XFILLER_4_529 VPWR VGND sg13g2_decap_8
XFILLER_0_735 VPWR VGND sg13g2_decap_8
XFILLER_48_728 VPWR VGND sg13g2_decap_8
XFILLER_47_238 VPWR VGND sg13g2_decap_8
XFILLER_46_21 VPWR VGND sg13g2_decap_8
XFILLER_29_942 VPWR VGND sg13g2_decap_8
XFILLER_44_901 VPWR VGND sg13g2_decap_8
XFILLER_28_463 VPWR VGND sg13g2_decap_8
XFILLER_46_98 VPWR VGND sg13g2_decap_8
XFILLER_43_411 VPWR VGND sg13g2_decap_8
XFILLER_15_102 VPWR VGND sg13g2_decap_8
XFILLER_16_636 VPWR VGND sg13g2_decap_8
XFILLER_44_978 VPWR VGND sg13g2_decap_8
XFILLER_31_617 VPWR VGND sg13g2_decap_8
XFILLER_43_488 VPWR VGND sg13g2_decap_8
XFILLER_8_802 VPWR VGND sg13g2_decap_8
XFILLER_23_190 VPWR VGND sg13g2_decap_8
XFILLER_30_138 VPWR VGND sg13g2_decap_8
XFILLER_7_301 VPWR VGND sg13g2_decap_8
XFILLER_12_886 VPWR VGND sg13g2_decap_8
XFILLER_8_879 VPWR VGND sg13g2_decap_8
XFILLER_11_396 VPWR VGND sg13g2_decap_8
X_125_ net13 VGND VPWR mod1.qam16_mod.q_level\[3\] mod1.q_out_qam16\[3\] clknet_2_0__leaf_clk
+ sg13g2_dfrbpq_1
XFILLER_7_378 VPWR VGND sg13g2_decap_8
X_056_ VPWR _032_ net4 VGND sg13g2_inv_1
XFILLER_39_739 VPWR VGND sg13g2_decap_8
XFILLER_38_249 VPWR VGND sg13g2_decap_8
XFILLER_19_496 VPWR VGND sg13g2_decap_8
XFILLER_34_433 VPWR VGND sg13g2_decap_8
XFILLER_35_934 VPWR VGND sg13g2_decap_8
XFILLER_21_116 VPWR VGND sg13g2_decap_8
XFILLER_22_639 VPWR VGND sg13g2_decap_8
XFILLER_38_750 VPWR VGND sg13g2_decap_8
XFILLER_44_208 VPWR VGND sg13g2_decap_8
XFILLER_25_411 VPWR VGND sg13g2_decap_8
XFILLER_26_945 VPWR VGND sg13g2_decap_8
XFILLER_37_271 VPWR VGND sg13g2_decap_8
XFILLER_41_915 VPWR VGND sg13g2_decap_8
XFILLER_13_606 VPWR VGND sg13g2_decap_8
XFILLER_16_46 VPWR VGND sg13g2_decap_8
XFILLER_12_116 VPWR VGND sg13g2_decap_8
XFILLER_25_488 VPWR VGND sg13g2_decap_8
XFILLER_40_425 VPWR VGND sg13g2_decap_8
XFILLER_8_109 VPWR VGND sg13g2_decap_8
XFILLER_32_12 VPWR VGND sg13g2_decap_8
XFILLER_21_661 VPWR VGND sg13g2_decap_8
XFILLER_20_193 VPWR VGND sg13g2_decap_8
XFILLER_32_89 VPWR VGND sg13g2_decap_8
XFILLER_5_816 VPWR VGND sg13g2_decap_8
XFILLER_4_326 VPWR VGND sg13g2_decap_8
XFILLER_0_532 VPWR VGND sg13g2_decap_8
XFILLER_48_525 VPWR VGND sg13g2_decap_8
XFILLER_16_433 VPWR VGND sg13g2_decap_8
XFILLER_17_945 VPWR VGND sg13g2_decap_8
XFILLER_44_775 VPWR VGND sg13g2_decap_8
XFILLER_32_915 VPWR VGND sg13g2_decap_8
XFILLER_43_285 VPWR VGND sg13g2_decap_8
XFILLER_31_414 VPWR VGND sg13g2_decap_8
XFILLER_12_683 VPWR VGND sg13g2_decap_8
XFILLER_40_992 VPWR VGND sg13g2_decap_8
XFILLER_8_676 VPWR VGND sg13g2_decap_8
XFILLER_7_175 VPWR VGND sg13g2_decap_8
XFILLER_11_193 VPWR VGND sg13g2_decap_8
X_108_ VPWR _005_ _023_ VGND sg13g2_inv_1
XFILLER_4_893 VPWR VGND sg13g2_decap_8
XFILLER_39_536 VPWR VGND sg13g2_decap_8
XFILLER_35_731 VPWR VGND sg13g2_decap_8
XFILLER_34_252 VPWR VGND sg13g2_decap_8
XFILLER_22_436 VPWR VGND sg13g2_decap_8
XFILLER_31_981 VPWR VGND sg13g2_decap_8
XFILLER_1_329 VPWR VGND sg13g2_decap_8
XFILLER_27_56 VPWR VGND sg13g2_decap_8
XFILLER_26_742 VPWR VGND sg13g2_decap_8
XFILLER_41_712 VPWR VGND sg13g2_decap_8
XFILLER_13_403 VPWR VGND sg13g2_decap_8
XFILLER_14_948 VPWR VGND sg13g2_decap_8
XFILLER_40_200 VPWR VGND sg13g2_decap_8
XFILLER_43_33 VPWR VGND sg13g2_decap_8
XFILLER_41_789 VPWR VGND sg13g2_decap_8
XFILLER_40_299 VPWR VGND sg13g2_decap_8
XFILLER_5_613 VPWR VGND sg13g2_decap_8
XFILLER_4_123 VPWR VGND sg13g2_decap_8
XFILLER_49_812 VPWR VGND sg13g2_decap_8
XFILLER_1_896 VPWR VGND sg13g2_decap_8
XFILLER_48_322 VPWR VGND sg13g2_decap_8
XFILLER_49_889 VPWR VGND sg13g2_decap_8
XFILLER_48_399 VPWR VGND sg13g2_decap_8
XFILLER_1_1001 VPWR VGND sg13g2_decap_8
XFILLER_17_742 VPWR VGND sg13g2_decap_8
XFILLER_44_572 VPWR VGND sg13g2_decap_8
XFILLER_16_263 VPWR VGND sg13g2_decap_8
XFILLER_32_712 VPWR VGND sg13g2_decap_8
XFILLER_31_222 VPWR VGND sg13g2_decap_8
XFILLER_13_970 VPWR VGND sg13g2_decap_8
XFILLER_20_929 VPWR VGND sg13g2_decap_8
XFILLER_32_789 VPWR VGND sg13g2_decap_8
XFILLER_9_963 VPWR VGND sg13g2_decap_8
XFILLER_12_480 VPWR VGND sg13g2_decap_8
XFILLER_31_288 VPWR VGND sg13g2_decap_8
XFILLER_8_473 VPWR VGND sg13g2_decap_8
XFILLER_4_690 VPWR VGND sg13g2_decap_8
XFILLER_39_311 VPWR VGND sg13g2_decap_8
XFILLER_27_539 VPWR VGND sg13g2_decap_8
XFILLER_42_509 VPWR VGND sg13g2_decap_8
XFILLER_11_907 VPWR VGND sg13g2_decap_8
XFILLER_22_233 VPWR VGND sg13g2_decap_8
XFILLER_23_767 VPWR VGND sg13g2_decap_8
Xfanout15 rst_n net15 VPWR VGND sg13g2_buf_8
XFILLER_10_417 VPWR VGND sg13g2_decap_8
XFILLER_13_25 VPWR VGND sg13g2_decap_8
XFILLER_22_299 VPWR VGND sg13g2_decap_8
XFILLER_2_627 VPWR VGND sg13g2_decap_8
XFILLER_1_126 VPWR VGND sg13g2_decap_8
XFILLER_49_119 VPWR VGND sg13g2_decap_8
XFILLER_38_11 VPWR VGND sg13g2_decap_8
XFILLER_46_826 VPWR VGND sg13g2_decap_8
XFILLER_38_88 VPWR VGND sg13g2_decap_8
XFILLER_45_369 VPWR VGND sg13g2_decap_8
XFILLER_33_509 VPWR VGND sg13g2_decap_8
XFILLER_13_200 VPWR VGND sg13g2_decap_8
XFILLER_14_745 VPWR VGND sg13g2_decap_8
XFILLER_41_586 VPWR VGND sg13g2_decap_8
XFILLER_13_277 VPWR VGND sg13g2_decap_8
XFILLER_6_900 VPWR VGND sg13g2_decap_8
XFILLER_5_410 VPWR VGND sg13g2_decap_8
XFILLER_10_984 VPWR VGND sg13g2_decap_8
XFILLER_6_977 VPWR VGND sg13g2_decap_8
XFILLER_5_487 VPWR VGND sg13g2_decap_8
XFILLER_1_693 VPWR VGND sg13g2_decap_8
XFILLER_37_804 VPWR VGND sg13g2_decap_8
XFILLER_49_686 VPWR VGND sg13g2_decap_8
XFILLER_48_196 VPWR VGND sg13g2_decap_8
XFILLER_36_347 VPWR VGND sg13g2_decap_8
XFILLER_20_726 VPWR VGND sg13g2_decap_8
XFILLER_32_586 VPWR VGND sg13g2_decap_8
XFILLER_9_760 VPWR VGND sg13g2_decap_8
XFILLER_30_1017 VPWR VGND sg13g2_decap_8
XFILLER_8_270 VPWR VGND sg13g2_decap_8
XFILLER_30_1028 VPWR VGND sg13g2_fill_1
XFILLER_5_81 VPWR VGND sg13g2_decap_8
XFILLER_39_130 VPWR VGND sg13g2_decap_8
XFILLER_28_848 VPWR VGND sg13g2_decap_8
XFILLER_27_336 VPWR VGND sg13g2_decap_8
XFILLER_42_306 VPWR VGND sg13g2_decap_8
XFILLER_11_704 VPWR VGND sg13g2_decap_8
XFILLER_23_564 VPWR VGND sg13g2_decap_8
XFILLER_24_46 VPWR VGND sg13g2_decap_8
XFILLER_10_214 VPWR VGND sg13g2_decap_8
XFILLER_6_207 VPWR VGND sg13g2_decap_8
XFILLER_40_67 VPWR VGND sg13g2_decap_8
XFILLER_3_914 VPWR VGND sg13g2_decap_8
XFILLER_49_21 VPWR VGND sg13g2_decap_8
XFILLER_6_4 VPWR VGND sg13g2_decap_8
XFILLER_2_424 VPWR VGND sg13g2_decap_8
XFILLER_49_98 VPWR VGND sg13g2_decap_8
XFILLER_1_28 VPWR VGND sg13g2_decap_8
XFILLER_19_804 VPWR VGND sg13g2_decap_8
XFILLER_46_623 VPWR VGND sg13g2_decap_8
XFILLER_18_347 VPWR VGND sg13g2_decap_8
XFILLER_34_818 VPWR VGND sg13g2_decap_8
XFILLER_45_166 VPWR VGND sg13g2_decap_8
XFILLER_42_873 VPWR VGND sg13g2_decap_8
XFILLER_14_542 VPWR VGND sg13g2_decap_8
XFILLER_41_383 VPWR VGND sg13g2_decap_8
XFILLER_10_781 VPWR VGND sg13g2_decap_8
XFILLER_6_774 VPWR VGND sg13g2_decap_8
XFILLER_5_284 VPWR VGND sg13g2_decap_8
XFILLER_39_4 VPWR VGND sg13g2_decap_8
XFILLER_2_991 VPWR VGND sg13g2_decap_8
XFILLER_1_490 VPWR VGND sg13g2_decap_8
XFILLER_37_601 VPWR VGND sg13g2_decap_8
XFILLER_49_483 VPWR VGND sg13g2_decap_8
Xinput5 ui_in[5] net5 VPWR VGND sg13g2_buf_2
XFILLER_24_306 VPWR VGND sg13g2_decap_8
XFILLER_36_166 VPWR VGND sg13g2_decap_8
XFILLER_37_678 VPWR VGND sg13g2_decap_8
XFILLER_33_873 VPWR VGND sg13g2_decap_8
XFILLER_20_523 VPWR VGND sg13g2_decap_8
XFILLER_32_383 VPWR VGND sg13g2_decap_8
XFILLER_0_917 VPWR VGND sg13g2_decap_8
XFILLER_19_46 VPWR VGND sg13g2_decap_8
XFILLER_27_133 VPWR VGND sg13g2_decap_8
XFILLER_28_645 VPWR VGND sg13g2_decap_8
XFILLER_42_103 VPWR VGND sg13g2_decap_8
XFILLER_16_818 VPWR VGND sg13g2_decap_8
XFILLER_35_12 VPWR VGND sg13g2_decap_8
XFILLER_24_851 VPWR VGND sg13g2_decap_8
XFILLER_35_89 VPWR VGND sg13g2_decap_8
XFILLER_11_501 VPWR VGND sg13g2_decap_8
XFILLER_23_361 VPWR VGND sg13g2_decap_8
X_141_ net13 VGND VPWR _014_ mod1.q_out_qpsk\[2\] clknet_2_2__leaf_clk sg13g2_dfrbpq_1
XFILLER_11_578 VPWR VGND sg13g2_decap_8
XFILLER_13_1012 VPWR VGND sg13g2_decap_8
X_072_ _043_ net22 VPWR VGND sg13g2_inv_4
XFILLER_3_711 VPWR VGND sg13g2_decap_8
XFILLER_2_221 VPWR VGND sg13g2_decap_8
XFILLER_3_788 VPWR VGND sg13g2_decap_8
XFILLER_2_298 VPWR VGND sg13g2_decap_8
XFILLER_47_910 VPWR VGND sg13g2_decap_8
XFILLER_19_601 VPWR VGND sg13g2_decap_8
XFILLER_46_420 VPWR VGND sg13g2_decap_8
XFILLER_20_1027 VPWR VGND sg13g2_fill_2
XFILLER_47_987 VPWR VGND sg13g2_decap_8
XFILLER_18_144 VPWR VGND sg13g2_decap_8
XFILLER_19_678 VPWR VGND sg13g2_decap_8
XFILLER_34_615 VPWR VGND sg13g2_decap_8
XFILLER_46_497 VPWR VGND sg13g2_decap_8
XFILLER_15_840 VPWR VGND sg13g2_decap_8
XFILLER_33_103 VPWR VGND sg13g2_decap_8
XFILLER_33_147 VPWR VGND sg13g2_fill_1
XFILLER_42_670 VPWR VGND sg13g2_decap_8
XFILLER_30_821 VPWR VGND sg13g2_decap_8
XFILLER_30_898 VPWR VGND sg13g2_decap_8
XFILLER_6_571 VPWR VGND sg13g2_decap_8
XFILLER_2_60 VPWR VGND sg13g2_decap_8
XFILLER_38_932 VPWR VGND sg13g2_decap_8
XFILLER_49_280 VPWR VGND sg13g2_decap_8
XFILLER_37_475 VPWR VGND sg13g2_decap_8
XFILLER_24_158 VPWR VGND sg13g2_decap_8
XFILLER_36_1012 VPWR VGND sg13g2_decap_8
XFILLER_40_607 VPWR VGND sg13g2_decap_8
XFILLER_33_670 VPWR VGND sg13g2_decap_8
XFILLER_21_843 VPWR VGND sg13g2_decap_8
XFILLER_32_180 VPWR VGND sg13g2_decap_8
XFILLER_21_25 VPWR VGND sg13g2_decap_8
XFILLER_4_508 VPWR VGND sg13g2_decap_8
XFILLER_0_714 VPWR VGND sg13g2_decap_8
XFILLER_48_707 VPWR VGND sg13g2_decap_8
XFILLER_43_1027 VPWR VGND sg13g2_fill_2
XFILLER_47_217 VPWR VGND sg13g2_decap_8
XFILLER_29_921 VPWR VGND sg13g2_decap_8
XFILLER_28_442 VPWR VGND sg13g2_decap_8
XFILLER_46_77 VPWR VGND sg13g2_decap_8
XFILLER_16_615 VPWR VGND sg13g2_decap_8
XFILLER_29_998 VPWR VGND sg13g2_decap_8
XFILLER_44_957 VPWR VGND sg13g2_decap_8
XFILLER_43_467 VPWR VGND sg13g2_decap_8
XFILLER_15_158 VPWR VGND sg13g2_decap_8
XFILLER_30_117 VPWR VGND sg13g2_decap_8
XFILLER_12_865 VPWR VGND sg13g2_decap_8
XFILLER_11_375 VPWR VGND sg13g2_decap_8
XFILLER_8_858 VPWR VGND sg13g2_decap_8
XFILLER_7_357 VPWR VGND sg13g2_decap_8
XFILLER_7_49 VPWR VGND sg13g2_decap_8
X_124_ net13 VGND VPWR mod1.qam16_mod.q_level\[2\] mod1.q_out_qam16\[2\] clknet_2_0__leaf_clk
+ sg13g2_dfrbpq_1
X_055_ VPWR mod1.qam16_mod.q_level\[3\] net3 VGND sg13g2_inv_1
XFILLER_3_585 VPWR VGND sg13g2_decap_8
XFILLER_39_718 VPWR VGND sg13g2_decap_8
XFILLER_38_228 VPWR VGND sg13g2_decap_8
XFILLER_47_784 VPWR VGND sg13g2_decap_8
XFILLER_19_475 VPWR VGND sg13g2_decap_8
XFILLER_35_913 VPWR VGND sg13g2_decap_8
XFILLER_46_294 VPWR VGND sg13g2_decap_8
XFILLER_34_412 VPWR VGND sg13g2_decap_8
XFILLER_22_618 VPWR VGND sg13g2_decap_8
XFILLER_34_489 VPWR VGND sg13g2_decap_8
XFILLER_30_695 VPWR VGND sg13g2_decap_8
XFILLER_26_924 VPWR VGND sg13g2_decap_8
XFILLER_37_250 VPWR VGND sg13g2_decap_8
XFILLER_16_25 VPWR VGND sg13g2_decap_8
XFILLER_25_467 VPWR VGND sg13g2_decap_8
XFILLER_40_404 VPWR VGND sg13g2_decap_8
XFILLER_21_640 VPWR VGND sg13g2_decap_8
XFILLER_20_172 VPWR VGND sg13g2_decap_8
XFILLER_32_68 VPWR VGND sg13g2_decap_8
XFILLER_4_305 VPWR VGND sg13g2_decap_8
XFILLER_10_1026 VPWR VGND sg13g2_fill_2
XFILLER_0_511 VPWR VGND sg13g2_decap_8
XFILLER_48_504 VPWR VGND sg13g2_decap_8
XFILLER_0_588 VPWR VGND sg13g2_decap_8
XFILLER_16_412 VPWR VGND sg13g2_decap_8
XFILLER_17_924 VPWR VGND sg13g2_decap_8
XFILLER_28_272 VPWR VGND sg13g2_decap_8
XFILLER_29_795 VPWR VGND sg13g2_decap_8
XFILLER_44_754 VPWR VGND sg13g2_decap_8
XFILLER_43_264 VPWR VGND sg13g2_decap_8
XFILLER_16_489 VPWR VGND sg13g2_decap_8
XFILLER_12_662 VPWR VGND sg13g2_decap_8
XFILLER_40_971 VPWR VGND sg13g2_decap_8
XFILLER_8_655 VPWR VGND sg13g2_decap_8
XFILLER_11_172 VPWR VGND sg13g2_decap_8
XFILLER_7_154 VPWR VGND sg13g2_decap_8
X_107_ net20 net12 _023_ VPWR VGND sg13g2_and2_1
XFILLER_4_872 VPWR VGND sg13g2_decap_8
XFILLER_3_382 VPWR VGND sg13g2_decap_8
XFILLER_26_1022 VPWR VGND sg13g2_decap_8
XFILLER_21_4 VPWR VGND sg13g2_decap_8
XFILLER_39_515 VPWR VGND sg13g2_decap_8
XFILLER_47_581 VPWR VGND sg13g2_decap_8
XFILLER_19_283 VPWR VGND sg13g2_fill_1
XFILLER_35_710 VPWR VGND sg13g2_decap_8
XFILLER_34_231 VPWR VGND sg13g2_decap_8
XFILLER_22_415 VPWR VGND sg13g2_decap_8
XFILLER_23_949 VPWR VGND sg13g2_decap_8
XFILLER_35_787 VPWR VGND sg13g2_decap_8
XFILLER_31_960 VPWR VGND sg13g2_decap_8
XFILLER_30_492 VPWR VGND sg13g2_decap_8
XFILLER_8_81 VPWR VGND sg13g2_decap_8
XFILLER_2_809 VPWR VGND sg13g2_decap_8
XFILLER_1_308 VPWR VGND sg13g2_decap_8
XFILLER_27_35 VPWR VGND sg13g2_decap_8
XFILLER_26_721 VPWR VGND sg13g2_decap_8
XFILLER_43_12 VPWR VGND sg13g2_decap_8
XFILLER_14_927 VPWR VGND sg13g2_decap_8
XFILLER_26_798 VPWR VGND sg13g2_decap_8
XFILLER_41_768 VPWR VGND sg13g2_decap_8
XFILLER_13_459 VPWR VGND sg13g2_decap_8
XFILLER_25_297 VPWR VGND sg13g2_decap_8
XFILLER_43_89 VPWR VGND sg13g2_decap_8
XFILLER_22_982 VPWR VGND sg13g2_decap_8
XFILLER_4_102 VPWR VGND sg13g2_decap_8
XFILLER_49_1022 VPWR VGND sg13g2_decap_8
XFILLER_5_669 VPWR VGND sg13g2_decap_8
XFILLER_4_179 VPWR VGND sg13g2_decap_8
XFILLER_4_39 VPWR VGND sg13g2_decap_8
XFILLER_48_301 VPWR VGND sg13g2_decap_8
XFILLER_1_875 VPWR VGND sg13g2_decap_8
XFILLER_49_868 VPWR VGND sg13g2_decap_8
XFILLER_0_385 VPWR VGND sg13g2_decap_8
XFILLER_48_378 VPWR VGND sg13g2_decap_8
XFILLER_17_721 VPWR VGND sg13g2_decap_8
XFILLER_36_529 VPWR VGND sg13g2_decap_8
XFILLER_44_551 VPWR VGND sg13g2_decap_8
XFILLER_16_242 VPWR VGND sg13g2_decap_8
XFILLER_29_592 VPWR VGND sg13g2_decap_8
XFILLER_17_798 VPWR VGND sg13g2_decap_8
XFILLER_31_201 VPWR VGND sg13g2_decap_8
XFILLER_20_908 VPWR VGND sg13g2_decap_8
XFILLER_31_267 VPWR VGND sg13g2_decap_8
XFILLER_32_768 VPWR VGND sg13g2_decap_8
XFILLER_9_942 VPWR VGND sg13g2_decap_8
XFILLER_8_452 VPWR VGND sg13g2_decap_8
XFILLER_27_518 VPWR VGND sg13g2_decap_8
XFILLER_39_389 VPWR VGND sg13g2_decap_8
XFILLER_22_201 VPWR VGND sg13g2_decap_8
XFILLER_35_584 VPWR VGND sg13g2_decap_8
XFILLER_22_223 VPWR VGND sg13g2_fill_1
XFILLER_23_746 VPWR VGND sg13g2_decap_8
XFILLER_2_606 VPWR VGND sg13g2_decap_8
XFILLER_1_105 VPWR VGND sg13g2_decap_8
XFILLER_46_805 VPWR VGND sg13g2_decap_8
XFILLER_38_67 VPWR VGND sg13g2_decap_8
XFILLER_18_529 VPWR VGND sg13g2_decap_8
XFILLER_45_348 VPWR VGND sg13g2_decap_8
XFILLER_14_724 VPWR VGND sg13g2_decap_8
XFILLER_26_595 VPWR VGND sg13g2_decap_8
XFILLER_41_565 VPWR VGND sg13g2_decap_8
XFILLER_13_256 VPWR VGND sg13g2_decap_8
XFILLER_9_249 VPWR VGND sg13g2_decap_8
XFILLER_16_1021 VPWR VGND sg13g2_decap_8
XFILLER_10_963 VPWR VGND sg13g2_decap_8
XFILLER_6_956 VPWR VGND sg13g2_decap_8
XFILLER_5_466 VPWR VGND sg13g2_decap_8
XFILLER_1_672 VPWR VGND sg13g2_decap_8
XFILLER_49_665 VPWR VGND sg13g2_decap_8
XFILLER_0_182 VPWR VGND sg13g2_decap_8
XFILLER_48_175 VPWR VGND sg13g2_decap_8
XFILLER_36_326 VPWR VGND sg13g2_decap_8
XFILLER_17_595 VPWR VGND sg13g2_decap_8
XFILLER_20_705 VPWR VGND sg13g2_decap_8
XFILLER_32_565 VPWR VGND sg13g2_decap_8
XFILLER_5_60 VPWR VGND sg13g2_decap_8
XFILLER_8_1019 VPWR VGND sg13g2_decap_8
XFILLER_27_315 VPWR VGND sg13g2_decap_8
XFILLER_28_827 VPWR VGND sg13g2_decap_8
XFILLER_39_186 VPWR VGND sg13g2_decap_8
XFILLER_35_381 VPWR VGND sg13g2_decap_8
XFILLER_36_893 VPWR VGND sg13g2_decap_8
XFILLER_23_543 VPWR VGND sg13g2_decap_8
XFILLER_24_25 VPWR VGND sg13g2_decap_8
XFILLER_40_46 VPWR VGND sg13g2_decap_8
XFILLER_2_403 VPWR VGND sg13g2_decap_8
XFILLER_49_77 VPWR VGND sg13g2_decap_8
XFILLER_46_602 VPWR VGND sg13g2_decap_8
XFILLER_18_326 VPWR VGND sg13g2_decap_8
XFILLER_45_145 VPWR VGND sg13g2_decap_8
XFILLER_46_679 VPWR VGND sg13g2_decap_8
XFILLER_27_882 VPWR VGND sg13g2_decap_8
XFILLER_14_521 VPWR VGND sg13g2_decap_8
XFILLER_26_392 VPWR VGND sg13g2_decap_8
XFILLER_42_852 VPWR VGND sg13g2_decap_8
XFILLER_41_362 VPWR VGND sg13g2_decap_8
XFILLER_14_598 VPWR VGND sg13g2_decap_8
XFILLER_10_760 VPWR VGND sg13g2_decap_8
XFILLER_6_753 VPWR VGND sg13g2_decap_8
XFILLER_5_263 VPWR VGND sg13g2_decap_8
XFILLER_2_970 VPWR VGND sg13g2_decap_8
XFILLER_49_462 VPWR VGND sg13g2_decap_8
Xinput6 ui_in[6] net6 VPWR VGND sg13g2_buf_2
XFILLER_37_657 VPWR VGND sg13g2_decap_8
XFILLER_36_145 VPWR VGND sg13g2_decap_8
XFILLER_18_893 VPWR VGND sg13g2_decap_8
XFILLER_17_392 VPWR VGND sg13g2_decap_8
XFILLER_33_852 VPWR VGND sg13g2_decap_8
XFILLER_20_502 VPWR VGND sg13g2_decap_8
XFILLER_32_362 VPWR VGND sg13g2_decap_8
XFILLER_20_579 VPWR VGND sg13g2_decap_8
XFILLER_19_25 VPWR VGND sg13g2_decap_8
XFILLER_28_624 VPWR VGND sg13g2_decap_8
XFILLER_27_112 VPWR VGND sg13g2_decap_8
XFILLER_43_649 VPWR VGND sg13g2_decap_8
XFILLER_24_830 VPWR VGND sg13g2_decap_8
XFILLER_27_189 VPWR VGND sg13g2_decap_8
XFILLER_36_690 VPWR VGND sg13g2_decap_8
XFILLER_42_159 VPWR VGND sg13g2_decap_8
XFILLER_23_340 VPWR VGND sg13g2_decap_8
XFILLER_35_68 VPWR VGND sg13g2_decap_8
XFILLER_11_557 VPWR VGND sg13g2_decap_8
X_140_ net14 VGND VPWR _003_ Demo1.epsk_de1.bit_out\[2\] clknet_2_1__leaf_clk sg13g2_dfrbpq_1
XFILLER_7_539 VPWR VGND sg13g2_decap_8
X_071_ _043_ _041_ Demo1.epsk_de1.bit_out\[1\] net11 Demo1.qam16_bits\[1\] VPWR VGND
+ sg13g2_a22oi_1
XFILLER_2_200 VPWR VGND sg13g2_decap_8
XFILLER_3_767 VPWR VGND sg13g2_decap_8
XFILLER_2_277 VPWR VGND sg13g2_decap_8
XFILLER_47_966 VPWR VGND sg13g2_decap_8
XFILLER_18_123 VPWR VGND sg13g2_decap_8
XFILLER_19_657 VPWR VGND sg13g2_decap_8
XFILLER_20_1006 VPWR VGND sg13g2_decap_8
XFILLER_46_476 VPWR VGND sg13g2_decap_8
XFILLER_15_896 VPWR VGND sg13g2_decap_8
XFILLER_30_800 VPWR VGND sg13g2_decap_8
XFILLER_14_395 VPWR VGND sg13g2_decap_8
XFILLER_30_877 VPWR VGND sg13g2_decap_8
XFILLER_6_550 VPWR VGND sg13g2_decap_8
XFILLER_38_911 VPWR VGND sg13g2_decap_8
XFILLER_37_454 VPWR VGND sg13g2_decap_8
XFILLER_38_988 VPWR VGND sg13g2_decap_8
XFILLER_18_690 VPWR VGND sg13g2_decap_8
XFILLER_25_649 VPWR VGND sg13g2_decap_8
XFILLER_24_137 VPWR VGND sg13g2_decap_8
XFILLER_21_822 VPWR VGND sg13g2_decap_8
XFILLER_20_365 VPWR VGND sg13g2_decap_8
XFILLER_21_899 VPWR VGND sg13g2_decap_8
XFILLER_43_1006 VPWR VGND sg13g2_decap_8
XFILLER_29_900 VPWR VGND sg13g2_decap_8
XFILLER_46_56 VPWR VGND sg13g2_decap_8
XFILLER_29_977 VPWR VGND sg13g2_decap_8
XFILLER_44_936 VPWR VGND sg13g2_decap_8
XFILLER_28_498 VPWR VGND sg13g2_decap_8
XFILLER_43_446 VPWR VGND sg13g2_decap_8
XFILLER_15_137 VPWR VGND sg13g2_decap_8
XFILLER_12_844 VPWR VGND sg13g2_decap_8
XFILLER_8_837 VPWR VGND sg13g2_decap_8
XFILLER_7_28 VPWR VGND sg13g2_decap_8
XFILLER_11_354 VPWR VGND sg13g2_decap_8
XFILLER_7_336 VPWR VGND sg13g2_decap_8
X_123_ _014_ _040_ mod1.qam16_mod.i_level\[3\] _039_ _035_ VPWR VGND sg13g2_a22oi_1
XFILLER_3_564 VPWR VGND sg13g2_decap_8
XFILLER_11_81 VPWR VGND sg13g2_decap_8
XFILLER_38_207 VPWR VGND sg13g2_decap_8
XFILLER_47_763 VPWR VGND sg13g2_decap_8
XFILLER_19_454 VPWR VGND sg13g2_decap_8
XFILLER_46_273 VPWR VGND sg13g2_decap_8
XFILLER_34_468 VPWR VGND sg13g2_decap_8
XFILLER_35_969 VPWR VGND sg13g2_decap_8
XFILLER_15_693 VPWR VGND sg13g2_decap_8
XFILLER_30_674 VPWR VGND sg13g2_decap_8
XFILLER_29_229 VPWR VGND sg13g2_decap_8
XFILLER_26_903 VPWR VGND sg13g2_decap_8
XFILLER_38_785 VPWR VGND sg13g2_decap_8
XFILLER_25_446 VPWR VGND sg13g2_decap_8
XFILLER_32_47 VPWR VGND sg13g2_decap_8
XFILLER_20_151 VPWR VGND sg13g2_decap_8
XFILLER_21_696 VPWR VGND sg13g2_decap_8
XFILLER_10_1005 VPWR VGND sg13g2_decap_8
XFILLER_0_567 VPWR VGND sg13g2_decap_8
XFILLER_17_903 VPWR VGND sg13g2_decap_8
XFILLER_29_774 VPWR VGND sg13g2_decap_8
XFILLER_44_733 VPWR VGND sg13g2_decap_8
XFILLER_43_243 VPWR VGND sg13g2_decap_8
XFILLER_16_468 VPWR VGND sg13g2_decap_8
XFILLER_31_449 VPWR VGND sg13g2_decap_8
XFILLER_12_641 VPWR VGND sg13g2_decap_8
XFILLER_40_950 VPWR VGND sg13g2_decap_8
XFILLER_8_634 VPWR VGND sg13g2_decap_8
XFILLER_11_151 VPWR VGND sg13g2_decap_8
XFILLER_7_133 VPWR VGND sg13g2_decap_8
X_106_ _032_ net5 _019_ _010_ VPWR VGND sg13g2_nor3_1
XFILLER_4_851 VPWR VGND sg13g2_decap_8
XFILLER_3_361 VPWR VGND sg13g2_decap_8
XFILLER_26_1001 VPWR VGND sg13g2_decap_8
XFILLER_14_4 VPWR VGND sg13g2_decap_8
XFILLER_47_560 VPWR VGND sg13g2_decap_8
XFILLER_19_262 VPWR VGND sg13g2_decap_8
XFILLER_34_210 VPWR VGND sg13g2_decap_8
XFILLER_35_766 VPWR VGND sg13g2_decap_8
XFILLER_23_928 VPWR VGND sg13g2_decap_8
XFILLER_15_490 VPWR VGND sg13g2_decap_8
XFILLER_34_287 VPWR VGND sg13g2_decap_8
XFILLER_34_298 VPWR VGND sg13g2_fill_2
XFILLER_8_60 VPWR VGND sg13g2_decap_8
XFILLER_30_471 VPWR VGND sg13g2_decap_8
XFILLER_33_1027 VPWR VGND sg13g2_fill_2
XFILLER_27_14 VPWR VGND sg13g2_decap_8
XFILLER_26_700 VPWR VGND sg13g2_decap_8
XFILLER_38_582 VPWR VGND sg13g2_decap_8
XFILLER_14_906 VPWR VGND sg13g2_decap_8
XFILLER_25_210 VPWR VGND sg13g2_fill_2
XFILLER_25_276 VPWR VGND sg13g2_decap_8
XFILLER_26_777 VPWR VGND sg13g2_decap_8
XFILLER_41_747 VPWR VGND sg13g2_decap_8
XFILLER_13_438 VPWR VGND sg13g2_decap_8
XFILLER_43_68 VPWR VGND sg13g2_decap_8
XFILLER_22_961 VPWR VGND sg13g2_decap_8
XFILLER_40_257 VPWR VGND sg13g2_decap_8
XFILLER_21_493 VPWR VGND sg13g2_decap_8
XFILLER_5_648 VPWR VGND sg13g2_decap_8
XFILLER_49_1001 VPWR VGND sg13g2_decap_8
XFILLER_4_158 VPWR VGND sg13g2_decap_8
XFILLER_4_18 VPWR VGND sg13g2_decap_8
XFILLER_1_854 VPWR VGND sg13g2_decap_8
XFILLER_0_364 VPWR VGND sg13g2_decap_8
XFILLER_49_847 VPWR VGND sg13g2_decap_8
XFILLER_48_357 VPWR VGND sg13g2_decap_8
XFILLER_36_508 VPWR VGND sg13g2_decap_8
XFILLER_17_700 VPWR VGND sg13g2_decap_8
XFILLER_29_571 VPWR VGND sg13g2_decap_8
XFILLER_44_530 VPWR VGND sg13g2_decap_8
XFILLER_16_221 VPWR VGND sg13g2_decap_8
XFILLER_17_91 VPWR VGND sg13g2_decap_8
XFILLER_17_777 VPWR VGND sg13g2_decap_8
XFILLER_16_298 VPWR VGND sg13g2_decap_8
XFILLER_32_747 VPWR VGND sg13g2_decap_8
XFILLER_9_921 VPWR VGND sg13g2_decap_8
XFILLER_31_246 VPWR VGND sg13g2_decap_8
XFILLER_8_431 VPWR VGND sg13g2_decap_8
XFILLER_9_998 VPWR VGND sg13g2_decap_8
XFILLER_39_368 VPWR VGND sg13g2_decap_8
XFILLER_35_563 VPWR VGND sg13g2_decap_8
XFILLER_23_725 VPWR VGND sg13g2_decap_8
XFILLER_22_268 VPWR VGND sg13g2_decap_4
XFILLER_18_508 VPWR VGND sg13g2_decap_8
XFILLER_38_46 VPWR VGND sg13g2_decap_8
XFILLER_45_327 VPWR VGND sg13g2_decap_8
XFILLER_14_703 VPWR VGND sg13g2_decap_8
XFILLER_26_574 VPWR VGND sg13g2_decap_8
XFILLER_41_544 VPWR VGND sg13g2_decap_8
XFILLER_13_235 VPWR VGND sg13g2_decap_8
XFILLER_16_1000 VPWR VGND sg13g2_decap_8
XFILLER_9_228 VPWR VGND sg13g2_decap_8
XFILLER_10_942 VPWR VGND sg13g2_decap_8
XFILLER_6_935 VPWR VGND sg13g2_decap_8
XFILLER_5_445 VPWR VGND sg13g2_decap_8
XFILLER_1_651 VPWR VGND sg13g2_decap_8
XFILLER_0_161 VPWR VGND sg13g2_decap_8
XFILLER_49_644 VPWR VGND sg13g2_decap_8
XFILLER_23_1026 VPWR VGND sg13g2_fill_2
XFILLER_48_154 VPWR VGND sg13g2_decap_8
XFILLER_36_305 VPWR VGND sg13g2_decap_8
XFILLER_37_839 VPWR VGND sg13g2_decap_8
XFILLER_17_574 VPWR VGND sg13g2_decap_8
XFILLER_45_894 VPWR VGND sg13g2_decap_8
XFILLER_32_544 VPWR VGND sg13g2_decap_8
XFILLER_9_795 VPWR VGND sg13g2_decap_8
XFILLER_28_806 VPWR VGND sg13g2_decap_8
XFILLER_39_165 VPWR VGND sg13g2_decap_8
XFILLER_36_872 VPWR VGND sg13g2_decap_8
XFILLER_23_522 VPWR VGND sg13g2_decap_8
XFILLER_35_360 VPWR VGND sg13g2_decap_8
XFILLER_11_739 VPWR VGND sg13g2_decap_8
XFILLER_23_599 VPWR VGND sg13g2_decap_8
XFILLER_10_249 VPWR VGND sg13g2_decap_8
XFILLER_40_25 VPWR VGND sg13g2_decap_8
XFILLER_46_1015 VPWR VGND sg13g2_decap_8
XFILLER_3_949 VPWR VGND sg13g2_decap_8
XFILLER_2_459 VPWR VGND sg13g2_decap_8
XFILLER_49_56 VPWR VGND sg13g2_decap_8
XFILLER_18_305 VPWR VGND sg13g2_decap_8
XFILLER_19_839 VPWR VGND sg13g2_decap_8
XFILLER_46_658 VPWR VGND sg13g2_decap_8
XFILLER_45_124 VPWR VGND sg13g2_decap_8
XFILLER_27_861 VPWR VGND sg13g2_decap_8
XFILLER_42_831 VPWR VGND sg13g2_decap_8
XFILLER_14_500 VPWR VGND sg13g2_decap_8
XFILLER_26_371 VPWR VGND sg13g2_decap_8
XFILLER_33_319 VPWR VGND sg13g2_decap_8
XFILLER_41_341 VPWR VGND sg13g2_decap_8
XFILLER_14_577 VPWR VGND sg13g2_decap_8
XFILLER_14_81 VPWR VGND sg13g2_decap_8
XFILLER_6_732 VPWR VGND sg13g2_decap_8
XFILLER_5_242 VPWR VGND sg13g2_decap_8
XFILLER_46_7 VPWR VGND sg13g2_decap_8
XFILLER_49_441 VPWR VGND sg13g2_decap_8
Xinput7 ui_in[7] net7 VPWR VGND sg13g2_buf_2
XFILLER_36_124 VPWR VGND sg13g2_decap_8
XFILLER_37_636 VPWR VGND sg13g2_decap_8
XFILLER_18_872 VPWR VGND sg13g2_decap_8
XFILLER_45_691 VPWR VGND sg13g2_decap_8
XFILLER_17_371 VPWR VGND sg13g2_decap_8
XFILLER_33_831 VPWR VGND sg13g2_decap_8
XFILLER_32_341 VPWR VGND sg13g2_decap_8
XFILLER_20_558 VPWR VGND sg13g2_decap_8
XFILLER_9_592 VPWR VGND sg13g2_decap_8
XFILLER_10_39 VPWR VGND sg13g2_decap_8
XFILLER_28_603 VPWR VGND sg13g2_decap_8
XFILLER_27_168 VPWR VGND sg13g2_decap_8
XFILLER_43_628 VPWR VGND sg13g2_decap_8
XFILLER_35_47 VPWR VGND sg13g2_decap_8
XFILLER_42_138 VPWR VGND sg13g2_decap_8
XFILLER_24_886 VPWR VGND sg13g2_decap_8
XFILLER_11_536 VPWR VGND sg13g2_decap_8
XFILLER_23_396 VPWR VGND sg13g2_decap_8
X_070_ _042_ net21 VPWR VGND sg13g2_inv_4
XFILLER_7_518 VPWR VGND sg13g2_decap_8
XFILLER_3_746 VPWR VGND sg13g2_decap_8
XFILLER_2_256 VPWR VGND sg13g2_decap_8
XFILLER_47_945 VPWR VGND sg13g2_decap_8
XFILLER_18_102 VPWR VGND sg13g2_decap_8
XFILLER_19_636 VPWR VGND sg13g2_decap_8
XFILLER_46_455 VPWR VGND sg13g2_decap_8
XFILLER_18_179 VPWR VGND sg13g2_decap_8
XFILLER_33_138 VPWR VGND sg13g2_decap_8
XFILLER_14_374 VPWR VGND sg13g2_decap_8
XFILLER_15_875 VPWR VGND sg13g2_decap_8
XFILLER_30_856 VPWR VGND sg13g2_decap_8
XFILLER_41_193 VPWR VGND sg13g2_decap_8
XFILLER_2_95 VPWR VGND sg13g2_decap_8
XFILLER_37_433 VPWR VGND sg13g2_decap_8
XFILLER_38_967 VPWR VGND sg13g2_decap_8
XFILLER_24_116 VPWR VGND sg13g2_decap_8
XFILLER_25_628 VPWR VGND sg13g2_decap_8
XFILLER_21_801 VPWR VGND sg13g2_decap_8
XFILLER_20_333 VPWR VGND sg13g2_decap_8
XFILLER_20_344 VPWR VGND sg13g2_fill_1
XFILLER_21_878 VPWR VGND sg13g2_decap_8
XFILLER_0_749 VPWR VGND sg13g2_decap_8
XFILLER_28_400 VPWR VGND sg13g2_fill_1
XFILLER_29_956 VPWR VGND sg13g2_decap_8
XFILLER_46_35 VPWR VGND sg13g2_decap_8
XFILLER_44_915 VPWR VGND sg13g2_decap_8
XFILLER_43_425 VPWR VGND sg13g2_decap_8
XFILLER_15_116 VPWR VGND sg13g2_decap_8
XFILLER_28_477 VPWR VGND sg13g2_decap_8
XFILLER_12_823 VPWR VGND sg13g2_decap_8
XFILLER_24_683 VPWR VGND sg13g2_decap_8
XFILLER_8_816 VPWR VGND sg13g2_decap_8
XFILLER_7_315 VPWR VGND sg13g2_decap_8
XFILLER_11_333 VPWR VGND sg13g2_decap_8
X_122_ net2 net48 _039_ _013_ VPWR VGND sg13g2_mux2_1
XFILLER_11_60 VPWR VGND sg13g2_decap_8
XFILLER_3_543 VPWR VGND sg13g2_decap_8
XFILLER_4_1012 VPWR VGND sg13g2_decap_8
XFILLER_19_433 VPWR VGND sg13g2_decap_8
XFILLER_47_742 VPWR VGND sg13g2_decap_8
XFILLER_46_252 VPWR VGND sg13g2_decap_8
XFILLER_35_948 VPWR VGND sg13g2_decap_8
XFILLER_34_447 VPWR VGND sg13g2_decap_8
XFILLER_15_672 VPWR VGND sg13g2_decap_8
XFILLER_43_992 VPWR VGND sg13g2_decap_8
XFILLER_14_193 VPWR VGND sg13g2_decap_8
XFILLER_30_653 VPWR VGND sg13g2_decap_8
Xinput10 uio_in[2] net10 VPWR VGND sg13g2_buf_1
XFILLER_7_882 VPWR VGND sg13g2_decap_8
XFILLER_38_764 VPWR VGND sg13g2_decap_8
XFILLER_25_425 VPWR VGND sg13g2_decap_8
XFILLER_37_285 VPWR VGND sg13g2_decap_8
XFILLER_26_959 VPWR VGND sg13g2_decap_8
XFILLER_41_929 VPWR VGND sg13g2_decap_8
XFILLER_40_439 VPWR VGND sg13g2_decap_8
XFILLER_20_130 VPWR VGND sg13g2_decap_8
XFILLER_32_26 VPWR VGND sg13g2_decap_8
XFILLER_21_675 VPWR VGND sg13g2_decap_8
XFILLER_10_1028 VPWR VGND sg13g2_fill_1
XFILLER_0_546 VPWR VGND sg13g2_decap_8
XFILLER_48_539 VPWR VGND sg13g2_decap_8
XFILLER_29_753 VPWR VGND sg13g2_decap_8
XFILLER_44_712 VPWR VGND sg13g2_decap_8
XFILLER_43_222 VPWR VGND sg13g2_decap_8
XFILLER_16_447 VPWR VGND sg13g2_decap_8
XFILLER_17_959 VPWR VGND sg13g2_decap_8
XFILLER_44_789 VPWR VGND sg13g2_decap_8
XFILLER_32_929 VPWR VGND sg13g2_decap_8
XFILLER_43_299 VPWR VGND sg13g2_decap_8
XFILLER_12_620 VPWR VGND sg13g2_decap_8
XFILLER_24_480 VPWR VGND sg13g2_decap_8
XFILLER_25_992 VPWR VGND sg13g2_decap_8
XFILLER_31_428 VPWR VGND sg13g2_decap_8
XFILLER_8_613 VPWR VGND sg13g2_decap_8
XFILLER_11_130 VPWR VGND sg13g2_decap_8
XFILLER_7_112 VPWR VGND sg13g2_decap_8
XFILLER_12_697 VPWR VGND sg13g2_decap_8
X_105_ net5 _040_ _019_ _009_ VPWR VGND sg13g2_nor3_1
XFILLER_7_189 VPWR VGND sg13g2_decap_8
XFILLER_22_81 VPWR VGND sg13g2_decap_8
XFILLER_4_830 VPWR VGND sg13g2_decap_8
XFILLER_3_340 VPWR VGND sg13g2_decap_8
XFILLER_19_241 VPWR VGND sg13g2_decap_8
XFILLER_23_907 VPWR VGND sg13g2_decap_8
XFILLER_35_745 VPWR VGND sg13g2_decap_8
XFILLER_34_266 VPWR VGND sg13g2_decap_8
XFILLER_33_1006 VPWR VGND sg13g2_decap_8
XFILLER_30_450 VPWR VGND sg13g2_decap_8
XFILLER_31_995 VPWR VGND sg13g2_decap_8
XFILLER_45_509 VPWR VGND sg13g2_decap_8
XFILLER_38_561 VPWR VGND sg13g2_decap_8
XFILLER_26_756 VPWR VGND sg13g2_decap_8
XFILLER_25_255 VPWR VGND sg13g2_decap_8
XFILLER_43_47 VPWR VGND sg13g2_decap_8
XFILLER_41_726 VPWR VGND sg13g2_decap_8
XFILLER_13_417 VPWR VGND sg13g2_decap_8
XFILLER_40_214 VPWR VGND sg13g2_fill_2
XFILLER_22_940 VPWR VGND sg13g2_decap_8
XFILLER_21_472 VPWR VGND sg13g2_decap_8
XFILLER_5_627 VPWR VGND sg13g2_decap_8
XFILLER_4_137 VPWR VGND sg13g2_decap_8
XFILLER_1_833 VPWR VGND sg13g2_decap_8
XFILLER_0_343 VPWR VGND sg13g2_decap_8
XFILLER_49_826 VPWR VGND sg13g2_decap_8
XFILLER_48_336 VPWR VGND sg13g2_decap_8
XFILLER_1_1015 VPWR VGND sg13g2_decap_8
XFILLER_29_550 VPWR VGND sg13g2_decap_8
XFILLER_16_200 VPWR VGND sg13g2_decap_8
XFILLER_17_756 VPWR VGND sg13g2_decap_8
XFILLER_17_70 VPWR VGND sg13g2_decap_8
XFILLER_44_586 VPWR VGND sg13g2_decap_8
XFILLER_16_277 VPWR VGND sg13g2_decap_8
XFILLER_32_726 VPWR VGND sg13g2_decap_8
XFILLER_9_900 VPWR VGND sg13g2_decap_8
XFILLER_8_410 VPWR VGND sg13g2_decap_8
XFILLER_13_984 VPWR VGND sg13g2_decap_8
XFILLER_9_977 VPWR VGND sg13g2_decap_8
XFILLER_12_494 VPWR VGND sg13g2_decap_8
XFILLER_8_487 VPWR VGND sg13g2_decap_8
XFILLER_39_325 VPWR VGND sg13g2_decap_8
XFILLER_23_704 VPWR VGND sg13g2_decap_8
XFILLER_35_542 VPWR VGND sg13g2_decap_8
XFILLER_22_247 VPWR VGND sg13g2_decap_8
XFILLER_13_39 VPWR VGND sg13g2_decap_8
XFILLER_31_792 VPWR VGND sg13g2_decap_8
XFILLER_38_25 VPWR VGND sg13g2_decap_8
XFILLER_45_306 VPWR VGND sg13g2_decap_8
XFILLER_26_553 VPWR VGND sg13g2_decap_8
XFILLER_41_523 VPWR VGND sg13g2_decap_8
XFILLER_13_214 VPWR VGND sg13g2_decap_8
XFILLER_9_207 VPWR VGND sg13g2_decap_8
XFILLER_14_759 VPWR VGND sg13g2_decap_8
XFILLER_10_921 VPWR VGND sg13g2_decap_8
XFILLER_21_291 VPWR VGND sg13g2_decap_8
XFILLER_6_914 VPWR VGND sg13g2_decap_8
XFILLER_5_424 VPWR VGND sg13g2_decap_8
XFILLER_10_998 VPWR VGND sg13g2_decap_8
XFILLER_1_630 VPWR VGND sg13g2_decap_8
XFILLER_49_623 VPWR VGND sg13g2_decap_8
XFILLER_0_140 VPWR VGND sg13g2_decap_8
XFILLER_23_1005 VPWR VGND sg13g2_decap_8
XFILLER_48_133 VPWR VGND sg13g2_decap_8
XFILLER_37_818 VPWR VGND sg13g2_decap_8
XFILLER_45_873 VPWR VGND sg13g2_decap_8
XFILLER_17_553 VPWR VGND sg13g2_decap_8
XFILLER_44_383 VPWR VGND sg13g2_decap_8
XFILLER_32_523 VPWR VGND sg13g2_decap_8
XFILLER_13_781 VPWR VGND sg13g2_decap_8
XFILLER_9_774 VPWR VGND sg13g2_decap_8
XFILLER_12_291 VPWR VGND sg13g2_decap_8
XFILLER_8_284 VPWR VGND sg13g2_decap_8
XFILLER_5_991 VPWR VGND sg13g2_decap_8
XFILLER_5_95 VPWR VGND sg13g2_decap_8
XFILLER_39_144 VPWR VGND sg13g2_decap_8
XFILLER_36_851 VPWR VGND sg13g2_decap_8
XFILLER_39_1012 VPWR VGND sg13g2_decap_8
XFILLER_23_501 VPWR VGND sg13g2_decap_8
XFILLER_11_718 VPWR VGND sg13g2_decap_8
XFILLER_23_578 VPWR VGND sg13g2_decap_8
XFILLER_10_228 VPWR VGND sg13g2_decap_8
XFILLER_3_928 VPWR VGND sg13g2_decap_8
XFILLER_2_438 VPWR VGND sg13g2_decap_8
XFILLER_49_35 VPWR VGND sg13g2_decap_8
XFILLER_19_818 VPWR VGND sg13g2_decap_8
XFILLER_46_637 VPWR VGND sg13g2_decap_8
XFILLER_45_103 VPWR VGND sg13g2_decap_8
XFILLER_27_840 VPWR VGND sg13g2_decap_8
XFILLER_42_810 VPWR VGND sg13g2_decap_8
XFILLER_26_350 VPWR VGND sg13g2_decap_8
XFILLER_41_320 VPWR VGND sg13g2_decap_8
XFILLER_14_556 VPWR VGND sg13g2_decap_8
XFILLER_42_887 VPWR VGND sg13g2_decap_8
XFILLER_41_397 VPWR VGND sg13g2_decap_8
XFILLER_14_60 VPWR VGND sg13g2_decap_8
XFILLER_6_711 VPWR VGND sg13g2_decap_8
XFILLER_5_221 VPWR VGND sg13g2_decap_8
XFILLER_10_795 VPWR VGND sg13g2_decap_8
XFILLER_6_788 VPWR VGND sg13g2_decap_8
XFILLER_5_298 VPWR VGND sg13g2_decap_8
XFILLER_49_420 VPWR VGND sg13g2_decap_8
Xinput8 uio_in[0] net8 VPWR VGND sg13g2_buf_1
XFILLER_37_615 VPWR VGND sg13g2_decap_8
XFILLER_49_497 VPWR VGND sg13g2_decap_8
XFILLER_36_103 VPWR VGND sg13g2_decap_8
XFILLER_18_851 VPWR VGND sg13g2_decap_8
XFILLER_45_670 VPWR VGND sg13g2_decap_8
XFILLER_17_350 VPWR VGND sg13g2_decap_8
XFILLER_33_810 VPWR VGND sg13g2_decap_8
XFILLER_44_180 VPWR VGND sg13g2_decap_8
XFILLER_32_320 VPWR VGND sg13g2_decap_8
XFILLER_33_887 VPWR VGND sg13g2_decap_8
XFILLER_20_537 VPWR VGND sg13g2_decap_8
XFILLER_32_397 VPWR VGND sg13g2_decap_8
XFILLER_9_571 VPWR VGND sg13g2_decap_8
XFILLER_10_18 VPWR VGND sg13g2_decap_8
XFILLER_43_607 VPWR VGND sg13g2_decap_8
XFILLER_27_147 VPWR VGND sg13g2_decap_8
XFILLER_28_659 VPWR VGND sg13g2_decap_8
XFILLER_42_117 VPWR VGND sg13g2_decap_8
XFILLER_15_309 VPWR VGND sg13g2_fill_2
XFILLER_35_26 VPWR VGND sg13g2_decap_8
XFILLER_24_865 VPWR VGND sg13g2_decap_8
XFILLER_35_180 VPWR VGND sg13g2_fill_2
XFILLER_11_515 VPWR VGND sg13g2_decap_8
XFILLER_23_375 VPWR VGND sg13g2_decap_8
XFILLER_13_1026 VPWR VGND sg13g2_fill_2
XFILLER_3_725 VPWR VGND sg13g2_decap_8
XFILLER_4_4 VPWR VGND sg13g2_decap_8
XFILLER_2_235 VPWR VGND sg13g2_decap_8
XFILLER_47_924 VPWR VGND sg13g2_decap_8
XFILLER_19_615 VPWR VGND sg13g2_decap_8
XFILLER_46_434 VPWR VGND sg13g2_decap_8
XFILLER_18_158 VPWR VGND sg13g2_decap_8
XFILLER_33_117 VPWR VGND sg13g2_decap_8
XFILLER_34_629 VPWR VGND sg13g2_decap_8
XFILLER_15_854 VPWR VGND sg13g2_decap_8
XFILLER_14_353 VPWR VGND sg13g2_decap_8
XFILLER_25_81 VPWR VGND sg13g2_decap_8
XFILLER_42_684 VPWR VGND sg13g2_decap_8
XFILLER_30_835 VPWR VGND sg13g2_decap_8
XFILLER_41_172 VPWR VGND sg13g2_decap_8
XFILLER_10_592 VPWR VGND sg13g2_decap_8
XFILLER_6_585 VPWR VGND sg13g2_decap_8
XFILLER_44_5 VPWR VGND sg13g2_decap_8
XFILLER_2_74 VPWR VGND sg13g2_decap_8
XFILLER_37_412 VPWR VGND sg13g2_decap_8
XFILLER_38_946 VPWR VGND sg13g2_decap_8
XFILLER_49_294 VPWR VGND sg13g2_decap_8
XFILLER_25_607 VPWR VGND sg13g2_decap_8
XFILLER_37_489 VPWR VGND sg13g2_decap_8
XFILLER_36_1026 VPWR VGND sg13g2_fill_2
XFILLER_20_312 VPWR VGND sg13g2_decap_8
XFILLER_33_684 VPWR VGND sg13g2_decap_8
XFILLER_21_857 VPWR VGND sg13g2_decap_8
XFILLER_32_194 VPWR VGND sg13g2_decap_8
XFILLER_21_39 VPWR VGND sg13g2_decap_8
XFILLER_0_728 VPWR VGND sg13g2_decap_8
XFILLER_46_14 VPWR VGND sg13g2_decap_8
XFILLER_29_935 VPWR VGND sg13g2_decap_8
XFILLER_28_456 VPWR VGND sg13g2_decap_8
XFILLER_43_404 VPWR VGND sg13g2_decap_8
XFILLER_16_629 VPWR VGND sg13g2_decap_8
XFILLER_12_802 VPWR VGND sg13g2_decap_8
XFILLER_24_662 VPWR VGND sg13g2_decap_8
XFILLER_11_312 VPWR VGND sg13g2_decap_8
XFILLER_23_172 VPWR VGND sg13g2_fill_2
XFILLER_23_183 VPWR VGND sg13g2_decap_8
XFILLER_12_879 VPWR VGND sg13g2_decap_8
X_121_ _012_ _039_ net46 VPWR VGND sg13g2_nand2b_1
XFILLER_11_389 VPWR VGND sg13g2_decap_8
XFILLER_3_522 VPWR VGND sg13g2_decap_8
XFILLER_3_599 VPWR VGND sg13g2_decap_8
XFILLER_47_721 VPWR VGND sg13g2_decap_8
XFILLER_19_412 VPWR VGND sg13g2_decap_8
XFILLER_46_231 VPWR VGND sg13g2_decap_8
XFILLER_47_798 VPWR VGND sg13g2_decap_8
XFILLER_19_489 VPWR VGND sg13g2_decap_8
XFILLER_35_927 VPWR VGND sg13g2_decap_8
XFILLER_34_426 VPWR VGND sg13g2_decap_8
XFILLER_43_971 VPWR VGND sg13g2_decap_8
XFILLER_15_651 VPWR VGND sg13g2_decap_8
XFILLER_21_109 VPWR VGND sg13g2_decap_8
XFILLER_42_481 VPWR VGND sg13g2_decap_8
XFILLER_14_172 VPWR VGND sg13g2_decap_8
XFILLER_30_632 VPWR VGND sg13g2_decap_8
Xinput11 uio_in[3] net16 VPWR VGND sg13g2_buf_1
XFILLER_7_861 VPWR VGND sg13g2_decap_8
XFILLER_6_382 VPWR VGND sg13g2_decap_8
XFILLER_38_743 VPWR VGND sg13g2_decap_8
XFILLER_26_938 VPWR VGND sg13g2_decap_8
XFILLER_37_264 VPWR VGND sg13g2_decap_8
XFILLER_41_908 VPWR VGND sg13g2_decap_8
XFILLER_16_39 VPWR VGND sg13g2_decap_8
XFILLER_12_109 VPWR VGND sg13g2_decap_8
XFILLER_40_418 VPWR VGND sg13g2_decap_8
XFILLER_33_481 VPWR VGND sg13g2_decap_8
XFILLER_34_993 VPWR VGND sg13g2_decap_8
XFILLER_21_654 VPWR VGND sg13g2_decap_8
XFILLER_5_809 VPWR VGND sg13g2_decap_8
XFILLER_20_186 VPWR VGND sg13g2_decap_8
XFILLER_4_319 VPWR VGND sg13g2_decap_8
XFILLER_0_525 VPWR VGND sg13g2_decap_8
XFILLER_48_518 VPWR VGND sg13g2_decap_8
XFILLER_29_732 VPWR VGND sg13g2_decap_8
XFILLER_43_201 VPWR VGND sg13g2_decap_8
XFILLER_17_938 VPWR VGND sg13g2_decap_8
XFILLER_16_426 VPWR VGND sg13g2_decap_8
XFILLER_28_286 VPWR VGND sg13g2_decap_4
XFILLER_44_768 VPWR VGND sg13g2_decap_8
XFILLER_25_971 VPWR VGND sg13g2_decap_8
XFILLER_31_407 VPWR VGND sg13g2_decap_8
XFILLER_32_908 VPWR VGND sg13g2_decap_8
XFILLER_43_278 VPWR VGND sg13g2_decap_8
XFILLER_19_1021 VPWR VGND sg13g2_decap_8
XFILLER_12_676 VPWR VGND sg13g2_decap_8
XFILLER_40_985 VPWR VGND sg13g2_decap_8
XFILLER_8_669 VPWR VGND sg13g2_decap_8
XFILLER_11_186 VPWR VGND sg13g2_decap_8
XFILLER_22_60 VPWR VGND sg13g2_decap_8
X_104_ _022_ VPWR _008_ VGND _039_ _020_ sg13g2_o21ai_1
XFILLER_7_168 VPWR VGND sg13g2_decap_8
XFILLER_4_886 VPWR VGND sg13g2_decap_8
XFILLER_3_396 VPWR VGND sg13g2_decap_8
XFILLER_39_529 VPWR VGND sg13g2_decap_8
XFILLER_19_220 VPWR VGND sg13g2_decap_8
XFILLER_35_724 VPWR VGND sg13g2_decap_8
XFILLER_47_595 VPWR VGND sg13g2_decap_8
XFILLER_19_297 VPWR VGND sg13g2_decap_8
XFILLER_34_245 VPWR VGND sg13g2_decap_8
XFILLER_16_993 VPWR VGND sg13g2_decap_8
XFILLER_22_429 VPWR VGND sg13g2_decap_8
XFILLER_31_974 VPWR VGND sg13g2_decap_8
XFILLER_8_95 VPWR VGND sg13g2_decap_8
XFILLER_38_540 VPWR VGND sg13g2_decap_8
XFILLER_27_49 VPWR VGND sg13g2_decap_8
XFILLER_25_212 VPWR VGND sg13g2_fill_1
XFILLER_26_735 VPWR VGND sg13g2_decap_8
XFILLER_41_705 VPWR VGND sg13g2_decap_8
XFILLER_43_26 VPWR VGND sg13g2_decap_8
XFILLER_34_790 VPWR VGND sg13g2_decap_8
XFILLER_21_451 VPWR VGND sg13g2_decap_8
XFILLER_22_996 VPWR VGND sg13g2_decap_8
XFILLER_5_606 VPWR VGND sg13g2_decap_8
XFILLER_4_116 VPWR VGND sg13g2_decap_8
XFILLER_1_812 VPWR VGND sg13g2_decap_8
XFILLER_49_805 VPWR VGND sg13g2_decap_8
XFILLER_0_322 VPWR VGND sg13g2_decap_8
XFILLER_48_315 VPWR VGND sg13g2_decap_8
XFILLER_1_889 VPWR VGND sg13g2_decap_8
XFILLER_0_399 VPWR VGND sg13g2_decap_8
XFILLER_17_735 VPWR VGND sg13g2_decap_8
XFILLER_44_565 VPWR VGND sg13g2_decap_8
XFILLER_16_256 VPWR VGND sg13g2_decap_8
XFILLER_32_705 VPWR VGND sg13g2_decap_8
XFILLER_31_215 VPWR VGND sg13g2_decap_8
XFILLER_13_963 VPWR VGND sg13g2_decap_8
XFILLER_12_473 VPWR VGND sg13g2_decap_8
XFILLER_40_782 VPWR VGND sg13g2_decap_8
XFILLER_9_956 VPWR VGND sg13g2_decap_8
XFILLER_8_466 VPWR VGND sg13g2_decap_8
XFILLER_4_683 VPWR VGND sg13g2_decap_8
XFILLER_3_193 VPWR VGND sg13g2_decap_8
XFILLER_39_304 VPWR VGND sg13g2_decap_8
XFILLER_48_882 VPWR VGND sg13g2_decap_8
XFILLER_47_392 VPWR VGND sg13g2_decap_8
XFILLER_35_521 VPWR VGND sg13g2_decap_8
XFILLER_35_598 VPWR VGND sg13g2_decap_8
XFILLER_16_790 VPWR VGND sg13g2_decap_8
XFILLER_13_18 VPWR VGND sg13g2_decap_8
XFILLER_31_771 VPWR VGND sg13g2_decap_8
XFILLER_30_292 VPWR VGND sg13g2_fill_2
XFILLER_1_119 VPWR VGND sg13g2_decap_8
XFILLER_46_819 VPWR VGND sg13g2_decap_8
XFILLER_26_532 VPWR VGND sg13g2_decap_8
XFILLER_39_893 VPWR VGND sg13g2_decap_8
XFILLER_41_502 VPWR VGND sg13g2_decap_8
XFILLER_14_738 VPWR VGND sg13g2_decap_8
XFILLER_41_579 VPWR VGND sg13g2_decap_8
XFILLER_10_900 VPWR VGND sg13g2_decap_8
XFILLER_21_270 VPWR VGND sg13g2_decap_8
XFILLER_22_793 VPWR VGND sg13g2_decap_8
XFILLER_5_403 VPWR VGND sg13g2_decap_8
XFILLER_10_977 VPWR VGND sg13g2_decap_8
XFILLER_49_602 VPWR VGND sg13g2_decap_8
XFILLER_1_686 VPWR VGND sg13g2_decap_8
XFILLER_48_112 VPWR VGND sg13g2_decap_8
XFILLER_0_196 VPWR VGND sg13g2_decap_8
XFILLER_23_1028 VPWR VGND sg13g2_fill_1
XFILLER_49_679 VPWR VGND sg13g2_decap_8
XFILLER_48_189 VPWR VGND sg13g2_decap_8
XFILLER_28_81 VPWR VGND sg13g2_decap_8
XFILLER_45_852 VPWR VGND sg13g2_decap_8
XFILLER_17_532 VPWR VGND sg13g2_decap_8
XFILLER_44_362 VPWR VGND sg13g2_decap_8
XFILLER_32_502 VPWR VGND sg13g2_decap_8
XFILLER_13_760 VPWR VGND sg13g2_decap_8
XFILLER_20_719 VPWR VGND sg13g2_decap_8
XFILLER_32_579 VPWR VGND sg13g2_decap_8
XFILLER_9_753 VPWR VGND sg13g2_decap_8
XFILLER_12_270 VPWR VGND sg13g2_decap_8
XFILLER_8_263 VPWR VGND sg13g2_decap_8
XFILLER_5_970 VPWR VGND sg13g2_decap_8
XFILLER_5_74 VPWR VGND sg13g2_decap_8
XFILLER_4_480 VPWR VGND sg13g2_decap_8
XFILLER_39_123 VPWR VGND sg13g2_decap_8
XFILLER_27_329 VPWR VGND sg13g2_decap_8
XFILLER_36_830 VPWR VGND sg13g2_decap_8
XFILLER_23_557 VPWR VGND sg13g2_decap_8
XFILLER_24_39 VPWR VGND sg13g2_decap_8
XFILLER_35_395 VPWR VGND sg13g2_decap_8
XFILLER_10_207 VPWR VGND sg13g2_decap_8
XFILLER_3_907 VPWR VGND sg13g2_decap_8
XFILLER_2_417 VPWR VGND sg13g2_decap_8
XFILLER_49_14 VPWR VGND sg13g2_decap_8
XFILLER_46_616 VPWR VGND sg13g2_decap_8
XFILLER_39_690 VPWR VGND sg13g2_decap_8
XFILLER_45_159 VPWR VGND sg13g2_decap_8
XFILLER_27_896 VPWR VGND sg13g2_decap_8
XFILLER_42_866 VPWR VGND sg13g2_decap_8
XFILLER_14_535 VPWR VGND sg13g2_decap_8
XFILLER_41_376 VPWR VGND sg13g2_decap_8
XFILLER_22_590 VPWR VGND sg13g2_decap_8
XFILLER_5_200 VPWR VGND sg13g2_decap_8
XFILLER_10_774 VPWR VGND sg13g2_decap_8
XFILLER_6_767 VPWR VGND sg13g2_decap_8
XFILLER_5_277 VPWR VGND sg13g2_decap_8
XFILLER_30_82 VPWR VGND sg13g2_decap_8
XFILLER_2_984 VPWR VGND sg13g2_decap_8
XFILLER_7_1022 VPWR VGND sg13g2_decap_8
XFILLER_1_483 VPWR VGND sg13g2_decap_8
XFILLER_49_476 VPWR VGND sg13g2_decap_8
XFILLER_18_830 VPWR VGND sg13g2_decap_8
Xinput9 uio_in[1] net9 VPWR VGND sg13g2_buf_1
XFILLER_36_159 VPWR VGND sg13g2_decap_8
XFILLER_33_866 VPWR VGND sg13g2_decap_8
XFILLER_20_516 VPWR VGND sg13g2_decap_8
XFILLER_32_376 VPWR VGND sg13g2_decap_8
XFILLER_9_550 VPWR VGND sg13g2_decap_8
XFILLER_19_39 VPWR VGND sg13g2_decap_8
XFILLER_27_126 VPWR VGND sg13g2_decap_8
XFILLER_28_638 VPWR VGND sg13g2_decap_8
XFILLER_24_844 VPWR VGND sg13g2_decap_8
XFILLER_35_192 VPWR VGND sg13g2_decap_8
XFILLER_23_354 VPWR VGND sg13g2_decap_8
XFILLER_13_1005 VPWR VGND sg13g2_decap_8
XFILLER_3_704 VPWR VGND sg13g2_decap_8
XFILLER_2_214 VPWR VGND sg13g2_decap_8
XFILLER_47_903 VPWR VGND sg13g2_decap_8
XFILLER_46_413 VPWR VGND sg13g2_decap_8
XFILLER_18_137 VPWR VGND sg13g2_decap_8
XFILLER_34_608 VPWR VGND sg13g2_decap_8
XFILLER_15_833 VPWR VGND sg13g2_decap_8
XFILLER_27_693 VPWR VGND sg13g2_decap_8
XFILLER_42_663 VPWR VGND sg13g2_decap_8
XFILLER_14_332 VPWR VGND sg13g2_decap_8
XFILLER_25_60 VPWR VGND sg13g2_decap_8
XFILLER_30_814 VPWR VGND sg13g2_decap_8
XFILLER_41_151 VPWR VGND sg13g2_decap_8
XFILLER_10_571 VPWR VGND sg13g2_decap_8
XFILLER_41_81 VPWR VGND sg13g2_decap_8
XFILLER_6_564 VPWR VGND sg13g2_decap_8
XFILLER_29_1012 VPWR VGND sg13g2_decap_8
XFILLER_2_781 VPWR VGND sg13g2_decap_8
XFILLER_1_280 VPWR VGND sg13g2_decap_8
XFILLER_2_53 VPWR VGND sg13g2_decap_8
XFILLER_49_273 VPWR VGND sg13g2_decap_8
XFILLER_38_925 VPWR VGND sg13g2_decap_8
XFILLER_46_980 VPWR VGND sg13g2_decap_8
XFILLER_37_468 VPWR VGND sg13g2_decap_8
XFILLER_33_663 VPWR VGND sg13g2_decap_8
XFILLER_36_1005 VPWR VGND sg13g2_decap_8
XFILLER_21_836 VPWR VGND sg13g2_decap_8
XFILLER_32_173 VPWR VGND sg13g2_decap_8
XFILLER_21_18 VPWR VGND sg13g2_decap_8
XFILLER_0_707 VPWR VGND sg13g2_decap_8
XFILLER_29_914 VPWR VGND sg13g2_decap_8
XFILLER_28_435 VPWR VGND sg13g2_decap_8
XFILLER_16_608 VPWR VGND sg13g2_decap_8
XFILLER_24_641 VPWR VGND sg13g2_decap_8
XFILLER_23_151 VPWR VGND sg13g2_decap_8
XFILLER_12_858 VPWR VGND sg13g2_decap_8
X_120_ _030_ _031_ _002_ VPWR VGND sg13g2_and2_1
XFILLER_11_368 VPWR VGND sg13g2_decap_8
XFILLER_20_880 VPWR VGND sg13g2_decap_8
XFILLER_3_501 VPWR VGND sg13g2_decap_8
XFILLER_3_578 VPWR VGND sg13g2_decap_8
XFILLER_11_95 VPWR VGND sg13g2_decap_8
XFILLER_47_700 VPWR VGND sg13g2_decap_8
XFILLER_46_210 VPWR VGND sg13g2_decap_8
XFILLER_35_906 VPWR VGND sg13g2_decap_8
XFILLER_47_777 VPWR VGND sg13g2_decap_8
XFILLER_19_468 VPWR VGND sg13g2_decap_8
XFILLER_34_405 VPWR VGND sg13g2_decap_8
XFILLER_46_287 VPWR VGND sg13g2_decap_8
XFILLER_15_630 VPWR VGND sg13g2_decap_8
XFILLER_27_490 VPWR VGND sg13g2_decap_8
XFILLER_43_950 VPWR VGND sg13g2_decap_8
XFILLER_42_460 VPWR VGND sg13g2_decap_8
XFILLER_14_151 VPWR VGND sg13g2_decap_8
XFILLER_30_611 VPWR VGND sg13g2_decap_8
Xinput12 uio_in[4] net17 VPWR VGND sg13g2_buf_2
XFILLER_30_688 VPWR VGND sg13g2_decap_8
XFILLER_7_840 VPWR VGND sg13g2_decap_8
XFILLER_6_361 VPWR VGND sg13g2_decap_8
XFILLER_42_1020 VPWR VGND sg13g2_decap_8
XFILLER_38_722 VPWR VGND sg13g2_decap_8
XFILLER_26_917 VPWR VGND sg13g2_decap_8
XFILLER_37_243 VPWR VGND sg13g2_decap_8
XFILLER_38_799 VPWR VGND sg13g2_decap_8
XFILLER_16_18 VPWR VGND sg13g2_decap_8
XFILLER_34_972 VPWR VGND sg13g2_decap_8
XFILLER_33_460 VPWR VGND sg13g2_decap_8
XFILLER_21_633 VPWR VGND sg13g2_decap_8
XFILLER_20_165 VPWR VGND sg13g2_decap_8
XFILLER_10_1019 VPWR VGND sg13g2_decap_8
XFILLER_0_504 VPWR VGND sg13g2_decap_8
XFILLER_29_711 VPWR VGND sg13g2_decap_8
XFILLER_28_232 VPWR VGND sg13g2_decap_8
XFILLER_16_405 VPWR VGND sg13g2_decap_8
XFILLER_17_917 VPWR VGND sg13g2_decap_8
XFILLER_28_243 VPWR VGND sg13g2_fill_2
XFILLER_29_788 VPWR VGND sg13g2_decap_8
XFILLER_44_747 VPWR VGND sg13g2_decap_8
XFILLER_43_257 VPWR VGND sg13g2_decap_8
XFILLER_19_1000 VPWR VGND sg13g2_decap_8
XFILLER_25_950 VPWR VGND sg13g2_decap_8
XFILLER_12_655 VPWR VGND sg13g2_decap_8
XFILLER_40_964 VPWR VGND sg13g2_decap_8
XFILLER_11_165 VPWR VGND sg13g2_decap_8
XFILLER_8_648 VPWR VGND sg13g2_decap_8
XFILLER_7_147 VPWR VGND sg13g2_decap_8
X_103_ _022_ VPWR _007_ VGND net2 _039_ sg13g2_o21ai_1
XFILLER_4_865 VPWR VGND sg13g2_decap_8
XFILLER_3_375 VPWR VGND sg13g2_decap_8
XFILLER_26_1015 VPWR VGND sg13g2_decap_8
XFILLER_39_508 VPWR VGND sg13g2_decap_8
XFILLER_47_574 VPWR VGND sg13g2_decap_8
XFILLER_47_91 VPWR VGND sg13g2_decap_8
XFILLER_35_703 VPWR VGND sg13g2_decap_8
XFILLER_19_276 VPWR VGND sg13g2_decap_8
XFILLER_34_224 VPWR VGND sg13g2_decap_8
XFILLER_22_408 VPWR VGND sg13g2_decap_8
XFILLER_16_972 VPWR VGND sg13g2_decap_8
XFILLER_31_953 VPWR VGND sg13g2_decap_8
XFILLER_8_74 VPWR VGND sg13g2_decap_8
XFILLER_30_485 VPWR VGND sg13g2_decap_8
XFILLER_26_714 VPWR VGND sg13g2_decap_8
XFILLER_27_28 VPWR VGND sg13g2_decap_8
XFILLER_38_596 VPWR VGND sg13g2_decap_8
XFILLER_21_430 VPWR VGND sg13g2_decap_8
XFILLER_22_975 VPWR VGND sg13g2_decap_8
XFILLER_49_1015 VPWR VGND sg13g2_decap_8
XFILLER_0_301 VPWR VGND sg13g2_decap_8
XFILLER_1_868 VPWR VGND sg13g2_decap_8
XFILLER_0_378 VPWR VGND sg13g2_decap_8
XFILLER_17_714 VPWR VGND sg13g2_decap_8
XFILLER_29_585 VPWR VGND sg13g2_decap_8
XFILLER_44_544 VPWR VGND sg13g2_decap_8
XFILLER_16_235 VPWR VGND sg13g2_decap_8
XFILLER_13_942 VPWR VGND sg13g2_decap_8
XFILLER_9_935 VPWR VGND sg13g2_decap_8
XFILLER_12_452 VPWR VGND sg13g2_decap_8
XFILLER_40_761 VPWR VGND sg13g2_decap_8
XFILLER_8_445 VPWR VGND sg13g2_decap_8
XFILLER_33_82 VPWR VGND sg13g2_decap_8
XFILLER_4_662 VPWR VGND sg13g2_decap_8
XFILLER_3_172 VPWR VGND sg13g2_decap_8
XFILLER_12_4 VPWR VGND sg13g2_decap_8
Xhold1 mod1.i_out_qpsk\[1\] VPWR VGND net46 sg13g2_dlygate4sd3_1
XFILLER_48_861 VPWR VGND sg13g2_decap_8
XFILLER_47_371 VPWR VGND sg13g2_decap_8
XFILLER_35_500 VPWR VGND sg13g2_decap_8
XFILLER_23_739 VPWR VGND sg13g2_decap_8
XFILLER_35_577 VPWR VGND sg13g2_decap_8
XFILLER_31_750 VPWR VGND sg13g2_decap_8
XFILLER_30_271 VPWR VGND sg13g2_decap_8
XFILLER_39_872 VPWR VGND sg13g2_decap_8
XFILLER_26_511 VPWR VGND sg13g2_decap_8
XFILLER_38_393 VPWR VGND sg13g2_decap_8
XFILLER_14_717 VPWR VGND sg13g2_decap_8
XFILLER_26_588 VPWR VGND sg13g2_decap_8
XFILLER_41_558 VPWR VGND sg13g2_decap_8
XFILLER_13_249 VPWR VGND sg13g2_decap_8
XFILLER_16_1014 VPWR VGND sg13g2_decap_8
XFILLER_22_772 VPWR VGND sg13g2_decap_8
XFILLER_10_956 VPWR VGND sg13g2_decap_8
XFILLER_6_949 VPWR VGND sg13g2_decap_8
XFILLER_5_459 VPWR VGND sg13g2_decap_8
XFILLER_1_665 VPWR VGND sg13g2_decap_8
XFILLER_49_658 VPWR VGND sg13g2_decap_8
XFILLER_0_175 VPWR VGND sg13g2_decap_8
XFILLER_48_168 VPWR VGND sg13g2_decap_8
XFILLER_45_831 VPWR VGND sg13g2_decap_8
XFILLER_17_511 VPWR VGND sg13g2_decap_8
XFILLER_28_60 VPWR VGND sg13g2_decap_8
XFILLER_29_382 VPWR VGND sg13g2_decap_8
XFILLER_36_319 VPWR VGND sg13g2_decap_8
XFILLER_44_341 VPWR VGND sg13g2_decap_8
XFILLER_17_588 VPWR VGND sg13g2_decap_8
XFILLER_32_558 VPWR VGND sg13g2_decap_8
XFILLER_9_732 VPWR VGND sg13g2_decap_8
XFILLER_8_242 VPWR VGND sg13g2_decap_8
XFILLER_5_53 VPWR VGND sg13g2_decap_8
XFILLER_39_102 VPWR VGND sg13g2_decap_8
XFILLER_27_308 VPWR VGND sg13g2_decap_8
XFILLER_39_179 VPWR VGND sg13g2_decap_8
XFILLER_35_374 VPWR VGND sg13g2_decap_8
XFILLER_36_886 VPWR VGND sg13g2_decap_8
XFILLER_23_536 VPWR VGND sg13g2_decap_8
XFILLER_24_18 VPWR VGND sg13g2_decap_8
XFILLER_40_39 VPWR VGND sg13g2_decap_8
XFILLER_18_319 VPWR VGND sg13g2_decap_8
XFILLER_45_138 VPWR VGND sg13g2_decap_8
XFILLER_14_514 VPWR VGND sg13g2_decap_8
XFILLER_27_875 VPWR VGND sg13g2_decap_8
XFILLER_42_845 VPWR VGND sg13g2_decap_8
XFILLER_26_385 VPWR VGND sg13g2_decap_8
XFILLER_41_355 VPWR VGND sg13g2_decap_8
XFILLER_10_753 VPWR VGND sg13g2_decap_8
XFILLER_14_95 VPWR VGND sg13g2_decap_8
XFILLER_6_746 VPWR VGND sg13g2_decap_8
XFILLER_5_256 VPWR VGND sg13g2_decap_8
XFILLER_30_61 VPWR VGND sg13g2_decap_8
XFILLER_7_1001 VPWR VGND sg13g2_decap_8
XFILLER_2_963 VPWR VGND sg13g2_decap_8
XFILLER_1_462 VPWR VGND sg13g2_decap_8
XFILLER_49_455 VPWR VGND sg13g2_decap_8
XFILLER_39_81 VPWR VGND sg13g2_decap_8
XFILLER_36_138 VPWR VGND sg13g2_decap_8
XFILLER_18_886 VPWR VGND sg13g2_decap_8
XFILLER_17_385 VPWR VGND sg13g2_decap_8
XFILLER_33_845 VPWR VGND sg13g2_decap_8
XFILLER_32_355 VPWR VGND sg13g2_decap_8
XFILLER_19_18 VPWR VGND sg13g2_decap_8
XFILLER_27_105 VPWR VGND sg13g2_decap_8
XFILLER_28_617 VPWR VGND sg13g2_decap_8
XFILLER_24_823 VPWR VGND sg13g2_decap_8
XFILLER_36_683 VPWR VGND sg13g2_decap_8
XFILLER_23_333 VPWR VGND sg13g2_decap_8
XFILLER_13_1028 VPWR VGND sg13g2_fill_1
XFILLER_18_116 VPWR VGND sg13g2_decap_8
XFILLER_47_959 VPWR VGND sg13g2_decap_8
XFILLER_46_469 VPWR VGND sg13g2_decap_8
XFILLER_15_812 VPWR VGND sg13g2_decap_8
XFILLER_27_672 VPWR VGND sg13g2_decap_8
XFILLER_14_311 VPWR VGND sg13g2_decap_8
XFILLER_42_642 VPWR VGND sg13g2_decap_8
XFILLER_15_889 VPWR VGND sg13g2_decap_8
XFILLER_41_130 VPWR VGND sg13g2_decap_8
XFILLER_14_388 VPWR VGND sg13g2_decap_8
XFILLER_10_550 VPWR VGND sg13g2_decap_8
XFILLER_6_543 VPWR VGND sg13g2_decap_8
XFILLER_41_60 VPWR VGND sg13g2_decap_8
XFILLER_2_760 VPWR VGND sg13g2_decap_8
XFILLER_2_32 VPWR VGND sg13g2_decap_8
XFILLER_38_904 VPWR VGND sg13g2_decap_8
XFILLER_49_252 VPWR VGND sg13g2_decap_8
XFILLER_37_447 VPWR VGND sg13g2_decap_8
XFILLER_17_182 VPWR VGND sg13g2_decap_8
XFILLER_18_683 VPWR VGND sg13g2_decap_8
XFILLER_33_642 VPWR VGND sg13g2_decap_8
XFILLER_21_815 VPWR VGND sg13g2_decap_8
XFILLER_32_152 VPWR VGND sg13g2_decap_8
XFILLER_36_1028 VPWR VGND sg13g2_fill_1
XFILLER_20_358 VPWR VGND sg13g2_decap_8
XFILLER_46_49 VPWR VGND sg13g2_decap_8
XFILLER_44_929 VPWR VGND sg13g2_decap_8
XFILLER_43_439 VPWR VGND sg13g2_decap_8
XFILLER_24_620 VPWR VGND sg13g2_decap_8
XFILLER_36_480 VPWR VGND sg13g2_decap_8
XFILLER_23_130 VPWR VGND sg13g2_decap_8
XFILLER_12_837 VPWR VGND sg13g2_decap_8
XFILLER_23_174 VPWR VGND sg13g2_fill_1
XFILLER_24_697 VPWR VGND sg13g2_decap_8
XFILLER_11_347 VPWR VGND sg13g2_decap_8
XFILLER_7_329 VPWR VGND sg13g2_decap_8
XFILLER_11_74 VPWR VGND sg13g2_decap_8
XFILLER_3_557 VPWR VGND sg13g2_decap_8
XFILLER_47_756 VPWR VGND sg13g2_decap_8
XFILLER_4_1026 VPWR VGND sg13g2_fill_2
XFILLER_19_447 VPWR VGND sg13g2_decap_8
XFILLER_46_266 VPWR VGND sg13g2_decap_8
XFILLER_28_981 VPWR VGND sg13g2_decap_8
XFILLER_36_82 VPWR VGND sg13g2_decap_8
XFILLER_14_130 VPWR VGND sg13g2_decap_8
XFILLER_15_686 VPWR VGND sg13g2_decap_8
Xinput13 uio_in[5] net18 VPWR VGND sg13g2_buf_2
XFILLER_30_667 VPWR VGND sg13g2_decap_8
XFILLER_6_340 VPWR VGND sg13g2_decap_8
XFILLER_7_896 VPWR VGND sg13g2_decap_8
XFILLER_38_701 VPWR VGND sg13g2_decap_8
XFILLER_37_222 VPWR VGND sg13g2_decap_8
XFILLER_38_778 VPWR VGND sg13g2_decap_8
XFILLER_18_480 VPWR VGND sg13g2_decap_8
XFILLER_25_439 VPWR VGND sg13g2_decap_8
XFILLER_37_299 VPWR VGND sg13g2_decap_8
XFILLER_34_951 VPWR VGND sg13g2_decap_8
XFILLER_21_612 VPWR VGND sg13g2_decap_8
XFILLER_20_144 VPWR VGND sg13g2_decap_8
XFILLER_21_689 VPWR VGND sg13g2_decap_8
XFILLER_28_211 VPWR VGND sg13g2_decap_8
Xclkbuf_2_2__f_clk clknet_0_clk clknet_2_2__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_29_767 VPWR VGND sg13g2_decap_8
XFILLER_44_726 VPWR VGND sg13g2_decap_8
XFILLER_43_236 VPWR VGND sg13g2_decap_8
XFILLER_12_634 VPWR VGND sg13g2_decap_8
XFILLER_24_494 VPWR VGND sg13g2_decap_8
XFILLER_40_943 VPWR VGND sg13g2_decap_8
XFILLER_8_627 VPWR VGND sg13g2_decap_8
XFILLER_11_144 VPWR VGND sg13g2_decap_8
XFILLER_7_126 VPWR VGND sg13g2_decap_8
X_102_ net4 mod1.qam16_mod.i_level\[3\] net3 _022_ VPWR VGND sg13g2_nand3_1
XFILLER_4_844 VPWR VGND sg13g2_decap_8
XFILLER_22_95 VPWR VGND sg13g2_decap_8
XFILLER_3_354 VPWR VGND sg13g2_decap_8
XFILLER_0_0 VPWR VGND sg13g2_decap_8
XFILLER_47_553 VPWR VGND sg13g2_decap_8
XFILLER_47_70 VPWR VGND sg13g2_decap_8
XFILLER_19_255 VPWR VGND sg13g2_decap_8
XFILLER_16_951 VPWR VGND sg13g2_decap_8
XFILLER_35_759 VPWR VGND sg13g2_decap_8
XFILLER_15_483 VPWR VGND sg13g2_decap_8
XFILLER_31_932 VPWR VGND sg13g2_decap_8
XFILLER_30_464 VPWR VGND sg13g2_decap_8
XFILLER_8_53 VPWR VGND sg13g2_decap_8
XFILLER_7_693 VPWR VGND sg13g2_decap_8
XFILLER_25_203 VPWR VGND sg13g2_decap_8
XFILLER_38_575 VPWR VGND sg13g2_decap_8
XFILLER_25_225 VPWR VGND sg13g2_decap_4
XFILLER_25_269 VPWR VGND sg13g2_decap_8
XFILLER_22_954 VPWR VGND sg13g2_decap_8
XFILLER_33_291 VPWR VGND sg13g2_decap_8
XFILLER_21_486 VPWR VGND sg13g2_decap_8
XFILLER_1_847 VPWR VGND sg13g2_decap_8
XFILLER_0_357 VPWR VGND sg13g2_decap_8
XFILLER_29_564 VPWR VGND sg13g2_decap_8
XFILLER_44_523 VPWR VGND sg13g2_decap_8
XFILLER_16_214 VPWR VGND sg13g2_decap_8
XFILLER_17_84 VPWR VGND sg13g2_decap_8
XFILLER_13_921 VPWR VGND sg13g2_decap_8
XFILLER_9_914 VPWR VGND sg13g2_decap_8
XFILLER_12_431 VPWR VGND sg13g2_decap_8
XFILLER_33_61 VPWR VGND sg13g2_decap_8
XFILLER_40_740 VPWR VGND sg13g2_decap_8
XFILLER_8_424 VPWR VGND sg13g2_decap_8
XFILLER_13_998 VPWR VGND sg13g2_decap_8
XFILLER_32_1020 VPWR VGND sg13g2_decap_8
XFILLER_4_641 VPWR VGND sg13g2_decap_8
XFILLER_3_151 VPWR VGND sg13g2_decap_8
Xhold2 mod1.q_out_qpsk\[2\] VPWR VGND net47 sg13g2_dlygate4sd3_1
XFILLER_48_840 VPWR VGND sg13g2_decap_8
XFILLER_47_350 VPWR VGND sg13g2_decap_8
XFILLER_35_556 VPWR VGND sg13g2_decap_8
XFILLER_23_718 VPWR VGND sg13g2_decap_8
XFILLER_30_250 VPWR VGND sg13g2_decap_8
XFILLER_8_991 VPWR VGND sg13g2_decap_8
XFILLER_7_490 VPWR VGND sg13g2_decap_8
XFILLER_38_39 VPWR VGND sg13g2_decap_8
XFILLER_39_851 VPWR VGND sg13g2_decap_8
XFILLER_38_361 VPWR VGND sg13g2_decap_8
XFILLER_38_372 VPWR VGND sg13g2_fill_1
XFILLER_26_567 VPWR VGND sg13g2_decap_8
XFILLER_41_537 VPWR VGND sg13g2_decap_8
XFILLER_13_228 VPWR VGND sg13g2_decap_8
XFILLER_22_751 VPWR VGND sg13g2_decap_8
XFILLER_10_935 VPWR VGND sg13g2_decap_8
XFILLER_6_928 VPWR VGND sg13g2_decap_8
XFILLER_5_438 VPWR VGND sg13g2_decap_8
XFILLER_1_644 VPWR VGND sg13g2_decap_8
XFILLER_0_154 VPWR VGND sg13g2_decap_8
XFILLER_49_637 VPWR VGND sg13g2_decap_8
XFILLER_23_1019 VPWR VGND sg13g2_decap_8
XFILLER_48_147 VPWR VGND sg13g2_decap_8
XFILLER_45_810 VPWR VGND sg13g2_decap_8
XFILLER_44_320 VPWR VGND sg13g2_decap_8
XFILLER_45_887 VPWR VGND sg13g2_decap_8
XFILLER_17_567 VPWR VGND sg13g2_decap_8
XFILLER_44_397 VPWR VGND sg13g2_decap_8
XFILLER_32_537 VPWR VGND sg13g2_decap_8
XFILLER_44_82 VPWR VGND sg13g2_decap_8
XFILLER_9_711 VPWR VGND sg13g2_decap_8
XFILLER_8_221 VPWR VGND sg13g2_decap_8
XFILLER_13_795 VPWR VGND sg13g2_decap_8
XFILLER_9_788 VPWR VGND sg13g2_decap_8
XFILLER_8_298 VPWR VGND sg13g2_decap_8
XFILLER_5_32 VPWR VGND sg13g2_decap_8
XFILLER_39_158 VPWR VGND sg13g2_decap_8
XFILLER_23_515 VPWR VGND sg13g2_decap_8
XFILLER_35_353 VPWR VGND sg13g2_decap_8
XFILLER_36_865 VPWR VGND sg13g2_decap_8
XFILLER_39_1026 VPWR VGND sg13g2_fill_2
XFILLER_40_18 VPWR VGND sg13g2_decap_8
XFILLER_46_1008 VPWR VGND sg13g2_decap_8
XFILLER_49_49 VPWR VGND sg13g2_decap_8
XFILLER_45_117 VPWR VGND sg13g2_decap_8
XFILLER_27_854 VPWR VGND sg13g2_decap_8
XFILLER_26_364 VPWR VGND sg13g2_decap_8
XFILLER_42_824 VPWR VGND sg13g2_decap_8
XFILLER_41_334 VPWR VGND sg13g2_decap_8
XFILLER_10_732 VPWR VGND sg13g2_decap_8
XFILLER_14_74 VPWR VGND sg13g2_decap_8
XFILLER_6_725 VPWR VGND sg13g2_decap_8
XFILLER_5_235 VPWR VGND sg13g2_decap_8
XFILLER_30_40 VPWR VGND sg13g2_decap_8
XFILLER_2_942 VPWR VGND sg13g2_decap_8
XFILLER_1_441 VPWR VGND sg13g2_decap_8
XFILLER_39_60 VPWR VGND sg13g2_decap_8
XFILLER_49_434 VPWR VGND sg13g2_decap_8
XFILLER_36_117 VPWR VGND sg13g2_decap_8
XFILLER_37_629 VPWR VGND sg13g2_decap_8
XFILLER_17_364 VPWR VGND sg13g2_decap_8
XFILLER_18_865 VPWR VGND sg13g2_decap_8
XFILLER_45_684 VPWR VGND sg13g2_decap_8
XFILLER_33_824 VPWR VGND sg13g2_decap_8
XFILLER_44_194 VPWR VGND sg13g2_decap_8
XFILLER_32_334 VPWR VGND sg13g2_decap_8
XFILLER_13_592 VPWR VGND sg13g2_decap_8
XFILLER_9_585 VPWR VGND sg13g2_decap_8
XFILLER_24_802 VPWR VGND sg13g2_decap_8
XFILLER_36_662 VPWR VGND sg13g2_decap_8
XFILLER_23_312 VPWR VGND sg13g2_decap_8
XFILLER_24_879 VPWR VGND sg13g2_decap_8
XFILLER_11_529 VPWR VGND sg13g2_decap_8
XFILLER_23_389 VPWR VGND sg13g2_decap_8
XFILLER_3_739 VPWR VGND sg13g2_decap_8
XFILLER_2_249 VPWR VGND sg13g2_decap_8
XFILLER_47_938 VPWR VGND sg13g2_decap_8
XFILLER_19_629 VPWR VGND sg13g2_decap_8
XFILLER_46_448 VPWR VGND sg13g2_decap_8
XFILLER_27_651 VPWR VGND sg13g2_decap_8
XFILLER_42_621 VPWR VGND sg13g2_decap_8
XFILLER_26_172 VPWR VGND sg13g2_decap_8
XFILLER_15_868 VPWR VGND sg13g2_decap_8
XFILLER_42_698 VPWR VGND sg13g2_decap_8
XFILLER_14_367 VPWR VGND sg13g2_decap_8
XFILLER_25_95 VPWR VGND sg13g2_decap_8
XFILLER_30_849 VPWR VGND sg13g2_decap_8
XFILLER_41_186 VPWR VGND sg13g2_decap_8
XFILLER_6_522 VPWR VGND sg13g2_decap_8
XFILLER_6_599 VPWR VGND sg13g2_decap_8
XFILLER_37_7 VPWR VGND sg13g2_decap_8
XFILLER_49_231 VPWR VGND sg13g2_decap_8
XFILLER_2_11 VPWR VGND sg13g2_decap_8
XFILLER_2_88 VPWR VGND sg13g2_decap_8
XFILLER_37_426 VPWR VGND sg13g2_decap_8
XFILLER_18_662 VPWR VGND sg13g2_decap_8
XFILLER_45_481 VPWR VGND sg13g2_decap_8
XFILLER_17_161 VPWR VGND sg13g2_decap_8
XFILLER_24_109 VPWR VGND sg13g2_decap_8
XFILLER_33_621 VPWR VGND sg13g2_decap_8
XFILLER_32_131 VPWR VGND sg13g2_decap_8
XFILLER_33_698 VPWR VGND sg13g2_decap_8
XFILLER_20_326 VPWR VGND sg13g2_decap_8
XFILLER_9_382 VPWR VGND sg13g2_decap_8
XFILLER_46_28 VPWR VGND sg13g2_decap_8
XFILLER_29_949 VPWR VGND sg13g2_decap_8
XFILLER_44_908 VPWR VGND sg13g2_decap_8
XFILLER_43_418 VPWR VGND sg13g2_decap_8
XFILLER_15_109 VPWR VGND sg13g2_decap_8
XFILLER_37_993 VPWR VGND sg13g2_decap_8
XFILLER_12_816 VPWR VGND sg13g2_decap_8
XFILLER_24_676 VPWR VGND sg13g2_decap_8
XFILLER_8_809 VPWR VGND sg13g2_decap_8
XFILLER_11_326 VPWR VGND sg13g2_decap_8
XFILLER_23_197 VPWR VGND sg13g2_decap_8
XFILLER_7_308 VPWR VGND sg13g2_decap_8
XFILLER_3_536 VPWR VGND sg13g2_decap_8
XFILLER_11_53 VPWR VGND sg13g2_decap_8
XFILLER_2_4 VPWR VGND sg13g2_decap_8
XFILLER_4_1005 VPWR VGND sg13g2_decap_8
XFILLER_47_735 VPWR VGND sg13g2_decap_8
XFILLER_19_426 VPWR VGND sg13g2_decap_8
XFILLER_46_245 VPWR VGND sg13g2_decap_8
XFILLER_28_960 VPWR VGND sg13g2_decap_8
XFILLER_36_61 VPWR VGND sg13g2_decap_8
XFILLER_43_985 VPWR VGND sg13g2_decap_8
XFILLER_15_665 VPWR VGND sg13g2_decap_8
XFILLER_42_495 VPWR VGND sg13g2_decap_8
XFILLER_14_186 VPWR VGND sg13g2_decap_8
XFILLER_30_646 VPWR VGND sg13g2_decap_8
Xinput14 uio_in[6] net19 VPWR VGND sg13g2_buf_2
XFILLER_11_893 VPWR VGND sg13g2_decap_8
XFILLER_7_875 VPWR VGND sg13g2_decap_8
XFILLER_6_396 VPWR VGND sg13g2_decap_8
XFILLER_42_5 VPWR VGND sg13g2_decap_8
XFILLER_37_201 VPWR VGND sg13g2_decap_8
XFILLER_38_757 VPWR VGND sg13g2_decap_8
XFILLER_19_993 VPWR VGND sg13g2_decap_8
XFILLER_25_418 VPWR VGND sg13g2_decap_8
XFILLER_37_278 VPWR VGND sg13g2_decap_8
XFILLER_34_930 VPWR VGND sg13g2_decap_8
XFILLER_20_123 VPWR VGND sg13g2_decap_8
XFILLER_32_19 VPWR VGND sg13g2_decap_8
XFILLER_33_495 VPWR VGND sg13g2_decap_8
XFILLER_21_668 VPWR VGND sg13g2_decap_8
XFILLER_0_539 VPWR VGND sg13g2_decap_8
XFILLER_29_746 VPWR VGND sg13g2_decap_8
XFILLER_44_705 VPWR VGND sg13g2_decap_8
XFILLER_43_215 VPWR VGND sg13g2_decap_8
XFILLER_37_790 VPWR VGND sg13g2_decap_8
XFILLER_12_613 VPWR VGND sg13g2_decap_8
XFILLER_25_985 VPWR VGND sg13g2_decap_8
XFILLER_40_922 VPWR VGND sg13g2_decap_8
XFILLER_11_123 VPWR VGND sg13g2_decap_8
XFILLER_24_473 VPWR VGND sg13g2_decap_8
XFILLER_8_606 VPWR VGND sg13g2_decap_8
XFILLER_7_105 VPWR VGND sg13g2_decap_8
X_101_ net5 _021_ _006_ VPWR VGND sg13g2_nor2_1
XFILLER_40_999 VPWR VGND sg13g2_decap_8
XFILLER_22_74 VPWR VGND sg13g2_decap_8
XFILLER_4_823 VPWR VGND sg13g2_decap_8
XFILLER_3_333 VPWR VGND sg13g2_decap_8
XFILLER_47_532 VPWR VGND sg13g2_decap_8
XFILLER_19_234 VPWR VGND sg13g2_decap_8
XFILLER_35_738 VPWR VGND sg13g2_decap_8
XFILLER_16_930 VPWR VGND sg13g2_decap_8
XFILLER_15_462 VPWR VGND sg13g2_decap_8
XFILLER_31_911 VPWR VGND sg13g2_decap_8
XFILLER_34_259 VPWR VGND sg13g2_decap_8
XFILLER_43_782 VPWR VGND sg13g2_decap_8
XFILLER_42_292 VPWR VGND sg13g2_decap_8
XFILLER_8_32 VPWR VGND sg13g2_decap_8
XFILLER_30_443 VPWR VGND sg13g2_decap_8
XFILLER_31_988 VPWR VGND sg13g2_decap_8
XFILLER_11_690 VPWR VGND sg13g2_decap_8
XFILLER_7_672 VPWR VGND sg13g2_decap_8
XFILLER_6_193 VPWR VGND sg13g2_decap_8
XFILLER_38_554 VPWR VGND sg13g2_decap_8
XFILLER_19_790 VPWR VGND sg13g2_decap_8
XFILLER_25_248 VPWR VGND sg13g2_decap_8
XFILLER_26_749 VPWR VGND sg13g2_decap_8
XFILLER_41_719 VPWR VGND sg13g2_decap_8
XFILLER_40_207 VPWR VGND sg13g2_decap_8
XFILLER_22_933 VPWR VGND sg13g2_decap_8
XFILLER_21_465 VPWR VGND sg13g2_decap_8
XFILLER_1_826 VPWR VGND sg13g2_decap_8
XFILLER_0_336 VPWR VGND sg13g2_decap_8
XFILLER_49_819 VPWR VGND sg13g2_decap_8
XFILLER_48_329 VPWR VGND sg13g2_decap_8
XFILLER_29_543 VPWR VGND sg13g2_decap_8
XFILLER_44_502 VPWR VGND sg13g2_decap_8
XFILLER_1_1008 VPWR VGND sg13g2_decap_8
XFILLER_17_63 VPWR VGND sg13g2_decap_8
XFILLER_17_749 VPWR VGND sg13g2_decap_8
XFILLER_44_579 VPWR VGND sg13g2_decap_8
XFILLER_13_900 VPWR VGND sg13g2_decap_8
XFILLER_32_719 VPWR VGND sg13g2_decap_8
XFILLER_12_410 VPWR VGND sg13g2_decap_8
XFILLER_25_782 VPWR VGND sg13g2_decap_8
XFILLER_8_403 VPWR VGND sg13g2_decap_8
XFILLER_13_977 VPWR VGND sg13g2_decap_8
XFILLER_24_292 VPWR VGND sg13g2_decap_8
XFILLER_33_40 VPWR VGND sg13g2_decap_8
XFILLER_12_487 VPWR VGND sg13g2_decap_8
XFILLER_40_796 VPWR VGND sg13g2_decap_8
XFILLER_4_620 VPWR VGND sg13g2_decap_8
XFILLER_3_130 VPWR VGND sg13g2_decap_8
XFILLER_4_697 VPWR VGND sg13g2_decap_8
Xhold3 mod1.i_out_qpsk\[2\] VPWR VGND net48 sg13g2_dlygate4sd3_1
XFILLER_39_318 VPWR VGND sg13g2_decap_8
XFILLER_48_896 VPWR VGND sg13g2_decap_8
XFILLER_35_535 VPWR VGND sg13g2_decap_8
XFILLER_22_218 VPWR VGND sg13g2_fill_2
XFILLER_31_785 VPWR VGND sg13g2_decap_8
XFILLER_8_970 VPWR VGND sg13g2_decap_8
XFILLER_38_18 VPWR VGND sg13g2_decap_8
XFILLER_39_830 VPWR VGND sg13g2_decap_8
XFILLER_38_340 VPWR VGND sg13g2_decap_8
XFILLER_26_546 VPWR VGND sg13g2_decap_8
XFILLER_41_516 VPWR VGND sg13g2_decap_8
XFILLER_13_207 VPWR VGND sg13g2_decap_8
XFILLER_22_730 VPWR VGND sg13g2_decap_8
XFILLER_10_914 VPWR VGND sg13g2_decap_8
XFILLER_6_907 VPWR VGND sg13g2_decap_8
XFILLER_21_284 VPWR VGND sg13g2_decap_8
XFILLER_5_417 VPWR VGND sg13g2_decap_8
XFILLER_1_623 VPWR VGND sg13g2_decap_8
XFILLER_49_616 VPWR VGND sg13g2_decap_8
XFILLER_0_133 VPWR VGND sg13g2_decap_8
XFILLER_48_126 VPWR VGND sg13g2_decap_8
XFILLER_17_546 VPWR VGND sg13g2_decap_8
XFILLER_28_95 VPWR VGND sg13g2_decap_8
XFILLER_45_866 VPWR VGND sg13g2_decap_8
XFILLER_44_376 VPWR VGND sg13g2_decap_8
XFILLER_44_61 VPWR VGND sg13g2_decap_8
XFILLER_32_516 VPWR VGND sg13g2_decap_8
XFILLER_8_200 VPWR VGND sg13g2_decap_8
XFILLER_13_774 VPWR VGND sg13g2_decap_8
XFILLER_9_767 VPWR VGND sg13g2_decap_8
XFILLER_12_284 VPWR VGND sg13g2_decap_8
XFILLER_40_593 VPWR VGND sg13g2_decap_8
XFILLER_8_277 VPWR VGND sg13g2_decap_8
XFILLER_5_11 VPWR VGND sg13g2_decap_8
XFILLER_5_984 VPWR VGND sg13g2_decap_8
XFILLER_5_88 VPWR VGND sg13g2_decap_8
XFILLER_4_494 VPWR VGND sg13g2_decap_8
XFILLER_39_137 VPWR VGND sg13g2_decap_8
XFILLER_48_693 VPWR VGND sg13g2_decap_8
XFILLER_35_332 VPWR VGND sg13g2_decap_8
XFILLER_36_844 VPWR VGND sg13g2_decap_8
XFILLER_39_1005 VPWR VGND sg13g2_decap_8
XFILLER_31_582 VPWR VGND sg13g2_decap_8
XFILLER_49_28 VPWR VGND sg13g2_decap_8
XFILLER_27_833 VPWR VGND sg13g2_decap_8
XFILLER_42_803 VPWR VGND sg13g2_decap_8
XFILLER_26_343 VPWR VGND sg13g2_decap_8
XFILLER_41_313 VPWR VGND sg13g2_decap_8
XFILLER_14_549 VPWR VGND sg13g2_decap_8
XFILLER_10_711 VPWR VGND sg13g2_decap_8
XFILLER_14_53 VPWR VGND sg13g2_decap_8
XFILLER_6_704 VPWR VGND sg13g2_decap_8
XFILLER_10_788 VPWR VGND sg13g2_decap_8
XFILLER_5_214 VPWR VGND sg13g2_decap_8
XFILLER_2_921 VPWR VGND sg13g2_decap_8
XFILLER_30_96 VPWR VGND sg13g2_decap_8
XFILLER_1_420 VPWR VGND sg13g2_decap_8
XFILLER_49_413 VPWR VGND sg13g2_decap_8
XFILLER_2_998 VPWR VGND sg13g2_decap_8
XFILLER_1_497 VPWR VGND sg13g2_decap_8
XFILLER_37_608 VPWR VGND sg13g2_decap_8
XFILLER_18_844 VPWR VGND sg13g2_decap_8
XFILLER_45_663 VPWR VGND sg13g2_decap_8
XFILLER_17_343 VPWR VGND sg13g2_decap_8
XFILLER_33_803 VPWR VGND sg13g2_decap_8
XFILLER_44_173 VPWR VGND sg13g2_decap_8
XFILLER_32_313 VPWR VGND sg13g2_decap_8
XFILLER_41_880 VPWR VGND sg13g2_decap_8
XFILLER_13_571 VPWR VGND sg13g2_decap_8
XFILLER_40_390 VPWR VGND sg13g2_decap_8
XFILLER_9_564 VPWR VGND sg13g2_decap_8
XFILLER_5_781 VPWR VGND sg13g2_decap_8
XFILLER_45_1020 VPWR VGND sg13g2_decap_8
XFILLER_4_291 VPWR VGND sg13g2_decap_8
XFILLER_49_980 VPWR VGND sg13g2_decap_8
XFILLER_48_490 VPWR VGND sg13g2_decap_8
XFILLER_35_19 VPWR VGND sg13g2_decap_8
XFILLER_36_641 VPWR VGND sg13g2_decap_8
XFILLER_35_173 VPWR VGND sg13g2_decap_8
XFILLER_24_858 VPWR VGND sg13g2_decap_8
XFILLER_11_508 VPWR VGND sg13g2_decap_8
XFILLER_23_368 VPWR VGND sg13g2_decap_8
XFILLER_32_880 VPWR VGND sg13g2_decap_8
XFILLER_13_1019 VPWR VGND sg13g2_decap_8
XFILLER_3_718 VPWR VGND sg13g2_decap_8
XFILLER_2_228 VPWR VGND sg13g2_decap_8
XFILLER_47_917 VPWR VGND sg13g2_decap_8
XFILLER_19_608 VPWR VGND sg13g2_decap_8
XFILLER_46_427 VPWR VGND sg13g2_decap_8
XFILLER_27_630 VPWR VGND sg13g2_decap_8
XFILLER_42_600 VPWR VGND sg13g2_decap_8
XFILLER_26_151 VPWR VGND sg13g2_decap_8
XFILLER_14_346 VPWR VGND sg13g2_decap_8
XFILLER_15_847 VPWR VGND sg13g2_decap_8
XFILLER_42_677 VPWR VGND sg13g2_decap_8
XFILLER_25_74 VPWR VGND sg13g2_decap_8
XFILLER_30_828 VPWR VGND sg13g2_decap_8
XFILLER_41_165 VPWR VGND sg13g2_decap_8
XFILLER_6_501 VPWR VGND sg13g2_decap_8
XFILLER_10_585 VPWR VGND sg13g2_decap_8
XFILLER_6_578 VPWR VGND sg13g2_decap_8
XFILLER_41_95 VPWR VGND sg13g2_decap_8
XFILLER_29_1026 VPWR VGND sg13g2_fill_2
XFILLER_49_210 VPWR VGND sg13g2_decap_8
XFILLER_2_795 VPWR VGND sg13g2_decap_8
XFILLER_1_294 VPWR VGND sg13g2_decap_8
XFILLER_2_67 VPWR VGND sg13g2_decap_8
XFILLER_37_405 VPWR VGND sg13g2_decap_8
XFILLER_38_939 VPWR VGND sg13g2_decap_8
XFILLER_49_287 VPWR VGND sg13g2_decap_8
XFILLER_18_641 VPWR VGND sg13g2_decap_8
XFILLER_46_994 VPWR VGND sg13g2_decap_8
XFILLER_45_460 VPWR VGND sg13g2_decap_8
XFILLER_17_140 VPWR VGND sg13g2_decap_8
XFILLER_33_600 VPWR VGND sg13g2_decap_8
XFILLER_32_110 VPWR VGND sg13g2_decap_8
XFILLER_20_305 VPWR VGND sg13g2_decap_8
XFILLER_33_677 VPWR VGND sg13g2_decap_8
XFILLER_36_1019 VPWR VGND sg13g2_decap_8
XFILLER_32_187 VPWR VGND sg13g2_decap_8
XFILLER_9_361 VPWR VGND sg13g2_decap_8
XFILLER_29_928 VPWR VGND sg13g2_decap_8
XFILLER_28_449 VPWR VGND sg13g2_decap_8
XFILLER_37_972 VPWR VGND sg13g2_decap_8
XFILLER_24_655 VPWR VGND sg13g2_decap_8
XFILLER_11_305 VPWR VGND sg13g2_decap_8
XFILLER_23_165 VPWR VGND sg13g2_decap_8
XFILLER_20_894 VPWR VGND sg13g2_decap_8
XFILLER_11_32 VPWR VGND sg13g2_decap_8
XFILLER_3_515 VPWR VGND sg13g2_decap_8
XFILLER_47_714 VPWR VGND sg13g2_decap_8
XFILLER_46_224 VPWR VGND sg13g2_decap_8
XFILLER_4_1028 VPWR VGND sg13g2_fill_1
XFILLER_34_419 VPWR VGND sg13g2_decap_8
XFILLER_36_40 VPWR VGND sg13g2_decap_8
XFILLER_15_644 VPWR VGND sg13g2_decap_8
XFILLER_43_964 VPWR VGND sg13g2_decap_8
XFILLER_42_474 VPWR VGND sg13g2_decap_8
XFILLER_14_165 VPWR VGND sg13g2_decap_8
XFILLER_30_625 VPWR VGND sg13g2_decap_8
Xinput15 uio_in[7] net20 VPWR VGND sg13g2_buf_2
XFILLER_11_872 VPWR VGND sg13g2_decap_8
XFILLER_10_382 VPWR VGND sg13g2_decap_8
XFILLER_7_854 VPWR VGND sg13g2_decap_8
XFILLER_6_375 VPWR VGND sg13g2_decap_8
XFILLER_2_592 VPWR VGND sg13g2_decap_8
XFILLER_35_5 VPWR VGND sg13g2_decap_8
XFILLER_28_4 VPWR VGND sg13g2_decap_8
XFILLER_38_736 VPWR VGND sg13g2_decap_8
XFILLER_37_257 VPWR VGND sg13g2_decap_8
XFILLER_19_972 VPWR VGND sg13g2_decap_8
XFILLER_46_791 VPWR VGND sg13g2_decap_8
XFILLER_34_986 VPWR VGND sg13g2_decap_8
XFILLER_20_102 VPWR VGND sg13g2_decap_8
XFILLER_21_647 VPWR VGND sg13g2_decap_8
XFILLER_33_474 VPWR VGND sg13g2_decap_8
XFILLER_20_179 VPWR VGND sg13g2_decap_8
XFILLER_0_518 VPWR VGND sg13g2_decap_8
XFILLER_29_725 VPWR VGND sg13g2_decap_8
XFILLER_16_419 VPWR VGND sg13g2_decap_8
XFILLER_28_279 VPWR VGND sg13g2_decap_8
XFILLER_19_1014 VPWR VGND sg13g2_decap_8
XFILLER_24_452 VPWR VGND sg13g2_decap_8
XFILLER_25_964 VPWR VGND sg13g2_decap_8
XFILLER_40_901 VPWR VGND sg13g2_decap_8
XFILLER_11_102 VPWR VGND sg13g2_decap_8
XFILLER_12_669 VPWR VGND sg13g2_decap_8
X_100_ _021_ net4 mod1.qam16_mod.q_level\[2\] VPWR VGND sg13g2_xnor2_1
XFILLER_40_978 VPWR VGND sg13g2_decap_8
XFILLER_11_179 VPWR VGND sg13g2_decap_8
XFILLER_4_802 VPWR VGND sg13g2_decap_8
XFILLER_20_691 VPWR VGND sg13g2_decap_8
XFILLER_22_53 VPWR VGND sg13g2_decap_8
XFILLER_3_312 VPWR VGND sg13g2_decap_8
XFILLER_4_879 VPWR VGND sg13g2_decap_8
XFILLER_3_389 VPWR VGND sg13g2_decap_8
XFILLER_47_511 VPWR VGND sg13g2_decap_8
XFILLER_19_213 VPWR VGND sg13g2_decap_8
XFILLER_47_588 VPWR VGND sg13g2_decap_8
XFILLER_35_717 VPWR VGND sg13g2_decap_8
XFILLER_34_238 VPWR VGND sg13g2_decap_8
XFILLER_43_761 VPWR VGND sg13g2_decap_8
XFILLER_15_441 VPWR VGND sg13g2_decap_8
XFILLER_16_986 VPWR VGND sg13g2_decap_8
XFILLER_42_271 VPWR VGND sg13g2_decap_8
XFILLER_30_422 VPWR VGND sg13g2_decap_8
XFILLER_8_11 VPWR VGND sg13g2_decap_8
XFILLER_31_967 VPWR VGND sg13g2_decap_8
XFILLER_8_88 VPWR VGND sg13g2_decap_8
XFILLER_7_651 VPWR VGND sg13g2_decap_8
XFILLER_30_499 VPWR VGND sg13g2_decap_8
XFILLER_6_172 VPWR VGND sg13g2_decap_8
XFILLER_38_533 VPWR VGND sg13g2_decap_8
XFILLER_26_728 VPWR VGND sg13g2_decap_8
XFILLER_43_19 VPWR VGND sg13g2_decap_8
XFILLER_22_912 VPWR VGND sg13g2_decap_8
XFILLER_34_783 VPWR VGND sg13g2_decap_8
XFILLER_21_444 VPWR VGND sg13g2_decap_8
XFILLER_22_989 VPWR VGND sg13g2_decap_8
XFILLER_4_109 VPWR VGND sg13g2_decap_8
XFILLER_1_805 VPWR VGND sg13g2_decap_8
XFILLER_0_315 VPWR VGND sg13g2_decap_8
XFILLER_48_308 VPWR VGND sg13g2_decap_8
XFILLER_29_522 VPWR VGND sg13g2_decap_8
XFILLER_17_728 VPWR VGND sg13g2_decap_8
XFILLER_17_42 VPWR VGND sg13g2_decap_8
XFILLER_29_599 VPWR VGND sg13g2_decap_8
XFILLER_44_558 VPWR VGND sg13g2_decap_8
XFILLER_16_249 VPWR VGND sg13g2_decap_8
XFILLER_25_761 VPWR VGND sg13g2_decap_8
XFILLER_31_208 VPWR VGND sg13g2_decap_8
XFILLER_24_271 VPWR VGND sg13g2_decap_8
XFILLER_13_956 VPWR VGND sg13g2_decap_8
XFILLER_9_949 VPWR VGND sg13g2_decap_8
XFILLER_12_466 VPWR VGND sg13g2_decap_8
XFILLER_40_775 VPWR VGND sg13g2_decap_8
XFILLER_8_459 VPWR VGND sg13g2_decap_8
XFILLER_33_96 VPWR VGND sg13g2_decap_8
XFILLER_4_676 VPWR VGND sg13g2_decap_8
XFILLER_3_186 VPWR VGND sg13g2_decap_8
XFILLER_0_882 VPWR VGND sg13g2_decap_8
XFILLER_48_875 VPWR VGND sg13g2_decap_8
XFILLER_35_514 VPWR VGND sg13g2_decap_8
XFILLER_47_385 VPWR VGND sg13g2_decap_8
XFILLER_16_783 VPWR VGND sg13g2_decap_8
XFILLER_22_208 VPWR VGND sg13g2_decap_8
XFILLER_31_764 VPWR VGND sg13g2_decap_8
XFILLER_30_285 VPWR VGND sg13g2_decap_8
XFILLER_39_886 VPWR VGND sg13g2_decap_8
XFILLER_26_525 VPWR VGND sg13g2_decap_8
XFILLER_34_580 VPWR VGND sg13g2_decap_8
XFILLER_16_1028 VPWR VGND sg13g2_fill_1
XFILLER_21_263 VPWR VGND sg13g2_decap_8
XFILLER_22_786 VPWR VGND sg13g2_decap_8
XFILLER_1_602 VPWR VGND sg13g2_decap_8
XFILLER_0_112 VPWR VGND sg13g2_decap_8
XFILLER_48_105 VPWR VGND sg13g2_decap_8
XFILLER_1_679 VPWR VGND sg13g2_decap_8
XFILLER_0_189 VPWR VGND sg13g2_decap_8
XFILLER_28_74 VPWR VGND sg13g2_decap_8
XFILLER_45_845 VPWR VGND sg13g2_decap_8
XFILLER_17_525 VPWR VGND sg13g2_decap_8
XFILLER_29_396 VPWR VGND sg13g2_decap_8
XFILLER_44_355 VPWR VGND sg13g2_decap_8
XFILLER_44_40 VPWR VGND sg13g2_decap_8
XFILLER_13_753 VPWR VGND sg13g2_decap_8
XFILLER_12_263 VPWR VGND sg13g2_decap_8
XFILLER_40_572 VPWR VGND sg13g2_decap_8
XFILLER_9_746 VPWR VGND sg13g2_decap_8
XFILLER_8_256 VPWR VGND sg13g2_decap_8
XFILLER_5_963 VPWR VGND sg13g2_decap_8
XFILLER_5_67 VPWR VGND sg13g2_decap_8
XFILLER_4_473 VPWR VGND sg13g2_decap_8
XFILLER_39_116 VPWR VGND sg13g2_decap_8
XFILLER_48_672 VPWR VGND sg13g2_decap_8
XFILLER_10_4 VPWR VGND sg13g2_decap_8
XFILLER_47_182 VPWR VGND sg13g2_decap_8
XFILLER_35_311 VPWR VGND sg13g2_decap_8
XFILLER_36_823 VPWR VGND sg13g2_decap_8
XFILLER_39_1028 VPWR VGND sg13g2_fill_1
XFILLER_35_388 VPWR VGND sg13g2_decap_8
XFILLER_16_580 VPWR VGND sg13g2_decap_8
XFILLER_31_561 VPWR VGND sg13g2_decap_8
XFILLER_46_609 VPWR VGND sg13g2_decap_8
XFILLER_22_1010 VPWR VGND sg13g2_decap_8
XFILLER_27_812 VPWR VGND sg13g2_decap_8
XFILLER_26_322 VPWR VGND sg13g2_decap_8
XFILLER_39_683 VPWR VGND sg13g2_decap_8
XFILLER_38_193 VPWR VGND sg13g2_decap_8
XFILLER_14_528 VPWR VGND sg13g2_decap_8
XFILLER_27_889 VPWR VGND sg13g2_decap_8
XFILLER_42_859 VPWR VGND sg13g2_decap_8
XFILLER_26_399 VPWR VGND sg13g2_decap_8
XFILLER_41_369 VPWR VGND sg13g2_decap_8
XFILLER_14_32 VPWR VGND sg13g2_decap_8
XFILLER_22_583 VPWR VGND sg13g2_decap_8
XFILLER_10_767 VPWR VGND sg13g2_decap_8
XFILLER_2_900 VPWR VGND sg13g2_decap_8
XFILLER_30_75 VPWR VGND sg13g2_decap_8
XFILLER_7_1015 VPWR VGND sg13g2_decap_8
XFILLER_2_977 VPWR VGND sg13g2_decap_8
XFILLER_1_476 VPWR VGND sg13g2_decap_8
XFILLER_49_469 VPWR VGND sg13g2_decap_8
XFILLER_39_95 VPWR VGND sg13g2_decap_8
XFILLER_17_322 VPWR VGND sg13g2_decap_8
XFILLER_18_823 VPWR VGND sg13g2_decap_8
XFILLER_45_642 VPWR VGND sg13g2_decap_8
XFILLER_29_182 VPWR VGND sg13g2_decap_8
XFILLER_29_193 VPWR VGND sg13g2_fill_2
XFILLER_44_152 VPWR VGND sg13g2_decap_8
XFILLER_17_399 VPWR VGND sg13g2_decap_8
XFILLER_33_859 VPWR VGND sg13g2_decap_8
XFILLER_13_550 VPWR VGND sg13g2_decap_8
XFILLER_20_509 VPWR VGND sg13g2_decap_8
XFILLER_32_369 VPWR VGND sg13g2_decap_8
XFILLER_9_543 VPWR VGND sg13g2_decap_8
XFILLER_5_760 VPWR VGND sg13g2_decap_8
XFILLER_4_270 VPWR VGND sg13g2_decap_8
XFILLER_27_119 VPWR VGND sg13g2_decap_8
XFILLER_36_620 VPWR VGND sg13g2_decap_8
XFILLER_24_837 VPWR VGND sg13g2_decap_8
XFILLER_35_152 VPWR VGND sg13g2_decap_8
XFILLER_36_697 VPWR VGND sg13g2_decap_8
XFILLER_23_347 VPWR VGND sg13g2_decap_8
XFILLER_2_207 VPWR VGND sg13g2_decap_8
XFILLER_46_406 VPWR VGND sg13g2_decap_8
XFILLER_39_480 VPWR VGND sg13g2_decap_8
XFILLER_26_130 VPWR VGND sg13g2_decap_8
XFILLER_15_826 VPWR VGND sg13g2_decap_8
XFILLER_27_686 VPWR VGND sg13g2_decap_8
XFILLER_42_656 VPWR VGND sg13g2_decap_8
XFILLER_14_325 VPWR VGND sg13g2_decap_8
XFILLER_25_53 VPWR VGND sg13g2_decap_8
XFILLER_30_807 VPWR VGND sg13g2_decap_8
XFILLER_41_144 VPWR VGND sg13g2_decap_8
XFILLER_10_564 VPWR VGND sg13g2_decap_8
XFILLER_41_74 VPWR VGND sg13g2_decap_8
XFILLER_6_557 VPWR VGND sg13g2_decap_8
XFILLER_29_1005 VPWR VGND sg13g2_decap_8
XFILLER_2_774 VPWR VGND sg13g2_decap_8
XFILLER_1_273 VPWR VGND sg13g2_decap_8
XFILLER_49_266 VPWR VGND sg13g2_decap_8
XFILLER_2_46 VPWR VGND sg13g2_decap_8
XFILLER_38_918 VPWR VGND sg13g2_decap_8
XFILLER_18_620 VPWR VGND sg13g2_decap_8
XFILLER_46_973 VPWR VGND sg13g2_decap_8
XFILLER_17_196 VPWR VGND sg13g2_decap_8
XFILLER_18_697 VPWR VGND sg13g2_decap_8
XFILLER_33_656 VPWR VGND sg13g2_decap_8
XFILLER_21_829 VPWR VGND sg13g2_decap_8
XFILLER_14_892 VPWR VGND sg13g2_decap_8
XFILLER_32_166 VPWR VGND sg13g2_decap_8
XFILLER_9_340 VPWR VGND sg13g2_decap_8
XFILLER_49_0 VPWR VGND sg13g2_decap_8
XFILLER_29_907 VPWR VGND sg13g2_decap_8
XFILLER_28_428 VPWR VGND sg13g2_decap_8
XFILLER_37_951 VPWR VGND sg13g2_decap_8
XFILLER_24_634 VPWR VGND sg13g2_decap_8
XFILLER_36_494 VPWR VGND sg13g2_decap_8
XFILLER_23_144 VPWR VGND sg13g2_decap_8
XFILLER_20_873 VPWR VGND sg13g2_decap_8
XFILLER_11_11 VPWR VGND sg13g2_decap_8
XFILLER_11_88 VPWR VGND sg13g2_decap_8
XFILLER_46_203 VPWR VGND sg13g2_decap_8
XFILLER_28_995 VPWR VGND sg13g2_decap_8
XFILLER_43_943 VPWR VGND sg13g2_decap_8
XFILLER_15_623 VPWR VGND sg13g2_decap_8
XFILLER_27_483 VPWR VGND sg13g2_decap_8
XFILLER_36_96 VPWR VGND sg13g2_decap_8
XFILLER_42_453 VPWR VGND sg13g2_decap_8
XFILLER_14_144 VPWR VGND sg13g2_decap_8
XFILLER_30_604 VPWR VGND sg13g2_decap_8
XFILLER_11_851 VPWR VGND sg13g2_decap_8
XFILLER_10_361 VPWR VGND sg13g2_decap_8
XFILLER_7_833 VPWR VGND sg13g2_decap_8
XFILLER_6_354 VPWR VGND sg13g2_decap_8
XFILLER_2_571 VPWR VGND sg13g2_decap_8
XFILLER_42_1013 VPWR VGND sg13g2_decap_8
XFILLER_38_715 VPWR VGND sg13g2_decap_8
XFILLER_19_951 VPWR VGND sg13g2_decap_8
XFILLER_37_236 VPWR VGND sg13g2_decap_8
XFILLER_46_770 VPWR VGND sg13g2_decap_8
XFILLER_18_494 VPWR VGND sg13g2_decap_8
XFILLER_33_453 VPWR VGND sg13g2_decap_8
XFILLER_34_965 VPWR VGND sg13g2_decap_8
XFILLER_21_626 VPWR VGND sg13g2_decap_8
XFILLER_20_158 VPWR VGND sg13g2_decap_8
XFILLER_29_704 VPWR VGND sg13g2_decap_8
XFILLER_28_225 VPWR VGND sg13g2_decap_8
XFILLER_25_943 VPWR VGND sg13g2_decap_8
XFILLER_24_431 VPWR VGND sg13g2_decap_8
XFILLER_12_648 VPWR VGND sg13g2_decap_8
XFILLER_40_957 VPWR VGND sg13g2_decap_8
XFILLER_11_158 VPWR VGND sg13g2_decap_8
XFILLER_20_670 VPWR VGND sg13g2_decap_8
XFILLER_22_32 VPWR VGND sg13g2_decap_8
XFILLER_4_858 VPWR VGND sg13g2_decap_8
XFILLER_3_368 VPWR VGND sg13g2_decap_8
XFILLER_26_1008 VPWR VGND sg13g2_decap_8
XFILLER_47_567 VPWR VGND sg13g2_decap_8
XFILLER_47_84 VPWR VGND sg13g2_decap_8
XFILLER_19_269 VPWR VGND sg13g2_decap_8
XFILLER_15_420 VPWR VGND sg13g2_decap_8
XFILLER_27_280 VPWR VGND sg13g2_decap_8
XFILLER_28_792 VPWR VGND sg13g2_decap_8
XFILLER_34_217 VPWR VGND sg13g2_decap_8
XFILLER_43_740 VPWR VGND sg13g2_decap_8
XFILLER_16_965 VPWR VGND sg13g2_decap_8
XFILLER_42_250 VPWR VGND sg13g2_decap_8
XFILLER_30_401 VPWR VGND sg13g2_decap_8
XFILLER_31_946 VPWR VGND sg13g2_decap_8
XFILLER_15_497 VPWR VGND sg13g2_decap_8
XFILLER_8_67 VPWR VGND sg13g2_decap_8
XFILLER_30_478 VPWR VGND sg13g2_decap_8
XFILLER_7_630 VPWR VGND sg13g2_decap_8
XFILLER_6_151 VPWR VGND sg13g2_decap_8
XFILLER_40_4 VPWR VGND sg13g2_decap_8
XFILLER_38_512 VPWR VGND sg13g2_decap_8
XFILLER_26_707 VPWR VGND sg13g2_decap_8
XFILLER_38_589 VPWR VGND sg13g2_decap_8
XFILLER_18_291 VPWR VGND sg13g2_decap_8
XFILLER_34_762 VPWR VGND sg13g2_decap_8
XFILLER_33_250 VPWR VGND sg13g2_decap_8
XFILLER_33_261 VPWR VGND sg13g2_fill_1
XFILLER_21_423 VPWR VGND sg13g2_decap_8
XFILLER_22_968 VPWR VGND sg13g2_decap_8
XFILLER_33_283 VPWR VGND sg13g2_fill_2
XFILLER_49_1008 VPWR VGND sg13g2_decap_8
XFILLER_29_501 VPWR VGND sg13g2_decap_8
XFILLER_17_21 VPWR VGND sg13g2_decap_8
XFILLER_17_707 VPWR VGND sg13g2_decap_8
XFILLER_29_578 VPWR VGND sg13g2_decap_8
XFILLER_44_537 VPWR VGND sg13g2_decap_8
XFILLER_16_228 VPWR VGND sg13g2_decap_8
XFILLER_17_98 VPWR VGND sg13g2_decap_8
XFILLER_25_740 VPWR VGND sg13g2_decap_8
XFILLER_13_935 VPWR VGND sg13g2_decap_8
XFILLER_24_250 VPWR VGND sg13g2_decap_8
XFILLER_12_445 VPWR VGND sg13g2_decap_8
XFILLER_40_754 VPWR VGND sg13g2_decap_8
XFILLER_9_928 VPWR VGND sg13g2_decap_8
XFILLER_33_75 VPWR VGND sg13g2_decap_8
XFILLER_8_438 VPWR VGND sg13g2_decap_8
XFILLER_21_990 VPWR VGND sg13g2_decap_8
XFILLER_4_655 VPWR VGND sg13g2_decap_8
XFILLER_3_165 VPWR VGND sg13g2_decap_8
XFILLER_0_861 VPWR VGND sg13g2_decap_8
XFILLER_48_854 VPWR VGND sg13g2_decap_8
XFILLER_47_364 VPWR VGND sg13g2_decap_8
XFILLER_15_261 VPWR VGND sg13g2_decap_8
XFILLER_16_762 VPWR VGND sg13g2_decap_8
XFILLER_31_743 VPWR VGND sg13g2_decap_8
XFILLER_30_264 VPWR VGND sg13g2_decap_8
XFILLER_30_297 VPWR VGND sg13g2_decap_8
XFILLER_26_504 VPWR VGND sg13g2_decap_8
XFILLER_39_865 VPWR VGND sg13g2_decap_8
XFILLER_38_386 VPWR VGND sg13g2_decap_8
XFILLER_16_1007 VPWR VGND sg13g2_decap_8
XFILLER_21_242 VPWR VGND sg13g2_decap_8
XFILLER_22_765 VPWR VGND sg13g2_decap_8
XFILLER_10_949 VPWR VGND sg13g2_decap_8
XFILLER_1_658 VPWR VGND sg13g2_decap_8
XFILLER_0_168 VPWR VGND sg13g2_decap_8
XFILLER_17_504 VPWR VGND sg13g2_decap_8
XFILLER_28_53 VPWR VGND sg13g2_decap_8
XFILLER_29_331 VPWR VGND sg13g2_decap_8
XFILLER_45_824 VPWR VGND sg13g2_decap_8
XFILLER_29_375 VPWR VGND sg13g2_decap_8
XFILLER_44_334 VPWR VGND sg13g2_decap_8
XFILLER_44_96 VPWR VGND sg13g2_decap_8
XFILLER_13_732 VPWR VGND sg13g2_decap_8
XFILLER_9_725 VPWR VGND sg13g2_decap_8
XFILLER_12_242 VPWR VGND sg13g2_decap_8
XFILLER_40_551 VPWR VGND sg13g2_decap_8
XFILLER_8_235 VPWR VGND sg13g2_decap_8
XFILLER_5_942 VPWR VGND sg13g2_decap_8
XFILLER_5_46 VPWR VGND sg13g2_decap_8
XFILLER_4_452 VPWR VGND sg13g2_decap_8
XFILLER_48_651 VPWR VGND sg13g2_decap_8
XFILLER_36_802 VPWR VGND sg13g2_decap_8
XFILLER_47_161 VPWR VGND sg13g2_decap_8
XFILLER_36_879 VPWR VGND sg13g2_decap_8
XFILLER_23_529 VPWR VGND sg13g2_decap_8
XFILLER_35_367 VPWR VGND sg13g2_decap_8
XFILLER_31_540 VPWR VGND sg13g2_decap_8
XFILLER_39_662 VPWR VGND sg13g2_decap_8
XFILLER_38_172 VPWR VGND sg13g2_decap_8
XFILLER_27_868 VPWR VGND sg13g2_decap_8
XFILLER_42_838 VPWR VGND sg13g2_decap_8
XFILLER_14_507 VPWR VGND sg13g2_decap_8
XFILLER_26_378 VPWR VGND sg13g2_decap_8
XFILLER_41_348 VPWR VGND sg13g2_decap_8
XFILLER_14_11 VPWR VGND sg13g2_decap_8
XFILLER_22_562 VPWR VGND sg13g2_decap_8
XFILLER_10_746 VPWR VGND sg13g2_decap_8
XFILLER_14_88 VPWR VGND sg13g2_decap_8
XFILLER_6_739 VPWR VGND sg13g2_decap_8
XFILLER_5_249 VPWR VGND sg13g2_decap_8
XFILLER_30_54 VPWR VGND sg13g2_decap_8
XFILLER_2_956 VPWR VGND sg13g2_decap_8
XFILLER_1_455 VPWR VGND sg13g2_decap_8
XFILLER_49_448 VPWR VGND sg13g2_decap_8
XFILLER_39_74 VPWR VGND sg13g2_decap_8
XFILLER_18_802 VPWR VGND sg13g2_decap_8
XFILLER_45_621 VPWR VGND sg13g2_decap_8
XFILLER_17_301 VPWR VGND sg13g2_decap_8
XFILLER_29_161 VPWR VGND sg13g2_decap_8
XFILLER_44_131 VPWR VGND sg13g2_decap_8
XFILLER_18_879 VPWR VGND sg13g2_decap_8
XFILLER_45_698 VPWR VGND sg13g2_decap_8
XFILLER_17_378 VPWR VGND sg13g2_decap_8
XFILLER_33_838 VPWR VGND sg13g2_decap_8
XFILLER_32_348 VPWR VGND sg13g2_decap_8
XFILLER_9_522 VPWR VGND sg13g2_decap_8
XFILLER_9_599 VPWR VGND sg13g2_decap_8
XFILLER_35_131 VPWR VGND sg13g2_decap_8
XFILLER_24_816 VPWR VGND sg13g2_decap_8
XFILLER_36_676 VPWR VGND sg13g2_decap_8
XFILLER_23_326 VPWR VGND sg13g2_decap_8
XFILLER_18_109 VPWR VGND sg13g2_decap_8
XFILLER_14_304 VPWR VGND sg13g2_decap_8
XFILLER_15_805 VPWR VGND sg13g2_decap_8
XFILLER_27_665 VPWR VGND sg13g2_decap_8
XFILLER_42_635 VPWR VGND sg13g2_decap_8
XFILLER_25_32 VPWR VGND sg13g2_decap_8
XFILLER_26_186 VPWR VGND sg13g2_decap_8
XFILLER_41_123 VPWR VGND sg13g2_decap_8
XFILLER_23_893 VPWR VGND sg13g2_decap_8
XFILLER_10_543 VPWR VGND sg13g2_decap_8
XFILLER_6_536 VPWR VGND sg13g2_decap_8
XFILLER_41_53 VPWR VGND sg13g2_decap_8
XFILLER_29_1028 VPWR VGND sg13g2_fill_1
XFILLER_2_753 VPWR VGND sg13g2_decap_8
XFILLER_1_252 VPWR VGND sg13g2_decap_8
XFILLER_2_25 VPWR VGND sg13g2_decap_8
XFILLER_49_245 VPWR VGND sg13g2_decap_8
XFILLER_46_952 VPWR VGND sg13g2_decap_8
XFILLER_18_676 VPWR VGND sg13g2_decap_8
XFILLER_45_495 VPWR VGND sg13g2_decap_8
XFILLER_17_175 VPWR VGND sg13g2_decap_8
XFILLER_33_635 VPWR VGND sg13g2_decap_8
XFILLER_21_808 VPWR VGND sg13g2_decap_8
XFILLER_32_145 VPWR VGND sg13g2_decap_8
XFILLER_14_871 VPWR VGND sg13g2_decap_8
XFILLER_9_396 VPWR VGND sg13g2_decap_8
XFILLER_37_930 VPWR VGND sg13g2_decap_8
XFILLER_24_613 VPWR VGND sg13g2_decap_8
XFILLER_36_473 VPWR VGND sg13g2_decap_8
XFILLER_23_123 VPWR VGND sg13g2_decap_8
XFILLER_20_852 VPWR VGND sg13g2_decap_8
XFILLER_11_67 VPWR VGND sg13g2_decap_8
XFILLER_4_1019 VPWR VGND sg13g2_decap_8
XFILLER_47_749 VPWR VGND sg13g2_decap_8
XFILLER_46_259 VPWR VGND sg13g2_decap_8
XFILLER_15_602 VPWR VGND sg13g2_decap_8
XFILLER_27_462 VPWR VGND sg13g2_decap_8
XFILLER_28_974 VPWR VGND sg13g2_decap_8
XFILLER_43_922 VPWR VGND sg13g2_decap_8
XFILLER_36_75 VPWR VGND sg13g2_decap_8
XFILLER_42_432 VPWR VGND sg13g2_decap_8
XFILLER_14_123 VPWR VGND sg13g2_decap_8
XFILLER_15_679 VPWR VGND sg13g2_decap_8
XFILLER_43_999 VPWR VGND sg13g2_decap_8
XFILLER_11_830 VPWR VGND sg13g2_decap_8
XFILLER_23_690 VPWR VGND sg13g2_decap_8
XFILLER_10_340 VPWR VGND sg13g2_decap_8
XFILLER_7_812 VPWR VGND sg13g2_decap_8
XFILLER_6_333 VPWR VGND sg13g2_decap_8
XFILLER_7_889 VPWR VGND sg13g2_decap_8
XFILLER_2_550 VPWR VGND sg13g2_decap_8
XFILLER_37_215 VPWR VGND sg13g2_decap_8
XFILLER_19_930 VPWR VGND sg13g2_decap_8
XFILLER_18_473 VPWR VGND sg13g2_decap_8
XFILLER_34_944 VPWR VGND sg13g2_decap_8
XFILLER_45_292 VPWR VGND sg13g2_decap_8
XFILLER_33_432 VPWR VGND sg13g2_decap_8
XFILLER_21_605 VPWR VGND sg13g2_decap_8
XFILLER_20_137 VPWR VGND sg13g2_decap_8
XFILLER_9_193 VPWR VGND sg13g2_decap_8
XFILLER_28_204 VPWR VGND sg13g2_decap_8
XFILLER_44_719 VPWR VGND sg13g2_decap_8
XFILLER_43_229 VPWR VGND sg13g2_decap_8
XFILLER_25_922 VPWR VGND sg13g2_decap_8
XFILLER_36_292 VPWR VGND sg13g2_fill_1
XFILLER_12_627 VPWR VGND sg13g2_decap_8
XFILLER_24_487 VPWR VGND sg13g2_decap_8
XFILLER_25_999 VPWR VGND sg13g2_decap_8
XFILLER_40_936 VPWR VGND sg13g2_decap_8
XFILLER_11_137 VPWR VGND sg13g2_decap_8
XFILLER_7_119 VPWR VGND sg13g2_decap_8
XFILLER_22_11 VPWR VGND sg13g2_decap_8
XFILLER_22_88 VPWR VGND sg13g2_decap_8
XFILLER_4_837 VPWR VGND sg13g2_decap_8
XFILLER_3_347 VPWR VGND sg13g2_decap_8
XFILLER_47_546 VPWR VGND sg13g2_decap_8
XFILLER_47_63 VPWR VGND sg13g2_decap_8
XFILLER_19_248 VPWR VGND sg13g2_decap_8
XFILLER_16_944 VPWR VGND sg13g2_decap_8
XFILLER_28_771 VPWR VGND sg13g2_decap_8
XFILLER_43_796 VPWR VGND sg13g2_decap_8
XFILLER_15_476 VPWR VGND sg13g2_decap_8
XFILLER_31_925 VPWR VGND sg13g2_decap_8
XFILLER_8_46 VPWR VGND sg13g2_decap_8
XFILLER_30_457 VPWR VGND sg13g2_decap_8
XFILLER_6_130 VPWR VGND sg13g2_decap_8
XFILLER_7_686 VPWR VGND sg13g2_decap_8
X_089_ _050_ _051_ _049_ net28 VPWR VGND _053_ sg13g2_nand4_1
XFILLER_38_568 VPWR VGND sg13g2_decap_8
XFILLER_18_270 VPWR VGND sg13g2_decap_8
XFILLER_25_218 VPWR VGND sg13g2_fill_2
XFILLER_25_229 VPWR VGND sg13g2_fill_2
XFILLER_34_741 VPWR VGND sg13g2_decap_8
XFILLER_21_402 VPWR VGND sg13g2_decap_8
XFILLER_22_947 VPWR VGND sg13g2_decap_8
XFILLER_21_479 VPWR VGND sg13g2_decap_8
XFILLER_25_1020 VPWR VGND sg13g2_decap_8
XFILLER_29_557 VPWR VGND sg13g2_decap_8
XFILLER_44_516 VPWR VGND sg13g2_decap_8
XFILLER_16_207 VPWR VGND sg13g2_decap_8
XFILLER_17_77 VPWR VGND sg13g2_decap_8
XFILLER_13_914 VPWR VGND sg13g2_decap_8
XFILLER_9_907 VPWR VGND sg13g2_decap_8
XFILLER_12_424 VPWR VGND sg13g2_decap_8
XFILLER_25_796 VPWR VGND sg13g2_decap_8
XFILLER_40_733 VPWR VGND sg13g2_decap_8
XFILLER_8_417 VPWR VGND sg13g2_decap_8
XFILLER_32_1013 VPWR VGND sg13g2_decap_8
XFILLER_33_54 VPWR VGND sg13g2_decap_8
XFILLER_4_634 VPWR VGND sg13g2_decap_8
XFILLER_3_144 VPWR VGND sg13g2_decap_8
XFILLER_0_840 VPWR VGND sg13g2_decap_8
XFILLER_48_833 VPWR VGND sg13g2_decap_8
XFILLER_47_343 VPWR VGND sg13g2_decap_8
XFILLER_16_741 VPWR VGND sg13g2_decap_8
XFILLER_35_549 VPWR VGND sg13g2_decap_8
XFILLER_15_240 VPWR VGND sg13g2_decap_8
XFILLER_43_593 VPWR VGND sg13g2_decap_8
XFILLER_15_295 VPWR VGND sg13g2_decap_8
XFILLER_31_722 VPWR VGND sg13g2_decap_8
XFILLER_30_243 VPWR VGND sg13g2_decap_8
XFILLER_12_991 VPWR VGND sg13g2_decap_8
XFILLER_31_799 VPWR VGND sg13g2_decap_8
XFILLER_8_984 VPWR VGND sg13g2_decap_8
XFILLER_7_483 VPWR VGND sg13g2_decap_8
XFILLER_39_844 VPWR VGND sg13g2_decap_8
XFILLER_38_354 VPWR VGND sg13g2_decap_8
XFILLER_0_1022 VPWR VGND sg13g2_decap_8
XFILLER_0_91 VPWR VGND sg13g2_decap_8
XFILLER_22_744 VPWR VGND sg13g2_decap_8
XFILLER_10_928 VPWR VGND sg13g2_decap_8
XFILLER_21_298 VPWR VGND sg13g2_decap_8
XFILLER_1_637 VPWR VGND sg13g2_decap_8
XFILLER_0_147 VPWR VGND sg13g2_decap_8
XFILLER_28_32 VPWR VGND sg13g2_decap_8
XFILLER_29_310 VPWR VGND sg13g2_decap_8
XFILLER_45_803 VPWR VGND sg13g2_decap_8
XFILLER_44_313 VPWR VGND sg13g2_decap_8
XFILLER_13_711 VPWR VGND sg13g2_decap_8
XFILLER_44_75 VPWR VGND sg13g2_decap_8
XFILLER_12_221 VPWR VGND sg13g2_decap_8
XFILLER_25_593 VPWR VGND sg13g2_decap_8
XFILLER_40_530 VPWR VGND sg13g2_decap_8
XFILLER_9_704 VPWR VGND sg13g2_decap_8
XFILLER_8_214 VPWR VGND sg13g2_decap_8
XFILLER_13_788 VPWR VGND sg13g2_decap_8
XFILLER_12_298 VPWR VGND sg13g2_decap_8
XFILLER_5_921 VPWR VGND sg13g2_decap_8
XFILLER_5_25 VPWR VGND sg13g2_decap_8
XFILLER_4_431 VPWR VGND sg13g2_decap_8
XFILLER_5_998 VPWR VGND sg13g2_decap_8
XFILLER_48_630 VPWR VGND sg13g2_decap_8
XFILLER_47_140 VPWR VGND sg13g2_decap_8
XFILLER_35_346 VPWR VGND sg13g2_decap_8
XFILLER_36_858 VPWR VGND sg13g2_decap_8
XFILLER_39_1019 VPWR VGND sg13g2_decap_8
XFILLER_23_508 VPWR VGND sg13g2_decap_8
XFILLER_44_880 VPWR VGND sg13g2_decap_8
XFILLER_43_390 VPWR VGND sg13g2_decap_8
XFILLER_31_596 VPWR VGND sg13g2_decap_8
XFILLER_8_781 VPWR VGND sg13g2_decap_8
XFILLER_7_280 VPWR VGND sg13g2_decap_8
XFILLER_39_641 VPWR VGND sg13g2_decap_8
XFILLER_38_151 VPWR VGND sg13g2_decap_8
XFILLER_27_847 VPWR VGND sg13g2_decap_8
XFILLER_42_817 VPWR VGND sg13g2_decap_8
XFILLER_26_357 VPWR VGND sg13g2_decap_8
XFILLER_41_327 VPWR VGND sg13g2_decap_8
XFILLER_22_541 VPWR VGND sg13g2_decap_8
XFILLER_10_725 VPWR VGND sg13g2_decap_8
XFILLER_14_67 VPWR VGND sg13g2_decap_8
XFILLER_6_718 VPWR VGND sg13g2_decap_8
XFILLER_5_228 VPWR VGND sg13g2_decap_8
XFILLER_30_33 VPWR VGND sg13g2_decap_8
XFILLER_2_935 VPWR VGND sg13g2_decap_8
XFILLER_1_434 VPWR VGND sg13g2_decap_8
XFILLER_49_427 VPWR VGND sg13g2_decap_8
XFILLER_39_53 VPWR VGND sg13g2_decap_8
XFILLER_45_600 VPWR VGND sg13g2_decap_8
XFILLER_29_140 VPWR VGND sg13g2_decap_8
XFILLER_44_110 VPWR VGND sg13g2_decap_8
XFILLER_18_858 VPWR VGND sg13g2_decap_8
XFILLER_45_677 VPWR VGND sg13g2_decap_8
XFILLER_17_357 VPWR VGND sg13g2_decap_8
XFILLER_33_817 VPWR VGND sg13g2_decap_8
XFILLER_44_187 VPWR VGND sg13g2_decap_8
XFILLER_32_327 VPWR VGND sg13g2_decap_8
XFILLER_9_501 VPWR VGND sg13g2_decap_8
XFILLER_41_894 VPWR VGND sg13g2_decap_8
XFILLER_13_585 VPWR VGND sg13g2_decap_8
XFILLER_9_578 VPWR VGND sg13g2_decap_8
XFILLER_5_795 VPWR VGND sg13g2_decap_8
XFILLER_49_994 VPWR VGND sg13g2_decap_8
XFILLER_35_110 VPWR VGND sg13g2_decap_8
XFILLER_36_655 VPWR VGND sg13g2_decap_8
XFILLER_23_305 VPWR VGND sg13g2_decap_8
XFILLER_32_894 VPWR VGND sg13g2_decap_8
XFILLER_31_393 VPWR VGND sg13g2_decap_8
XFILLER_27_644 VPWR VGND sg13g2_decap_8
XFILLER_25_11 VPWR VGND sg13g2_decap_8
XFILLER_42_614 VPWR VGND sg13g2_decap_8
XFILLER_26_165 VPWR VGND sg13g2_decap_8
XFILLER_41_102 VPWR VGND sg13g2_decap_8
XFILLER_25_88 VPWR VGND sg13g2_decap_8
XFILLER_23_872 VPWR VGND sg13g2_decap_8
XFILLER_41_179 VPWR VGND sg13g2_decap_8
XFILLER_10_522 VPWR VGND sg13g2_decap_8
XFILLER_41_32 VPWR VGND sg13g2_decap_8
XFILLER_6_515 VPWR VGND sg13g2_decap_8
XFILLER_10_599 VPWR VGND sg13g2_decap_8
XFILLER_2_732 VPWR VGND sg13g2_decap_8
XFILLER_1_231 VPWR VGND sg13g2_decap_8
XFILLER_49_224 VPWR VGND sg13g2_decap_8
XFILLER_37_419 VPWR VGND sg13g2_decap_8
XFILLER_46_931 VPWR VGND sg13g2_decap_8
XFILLER_17_154 VPWR VGND sg13g2_decap_8
XFILLER_18_655 VPWR VGND sg13g2_decap_8
XFILLER_45_474 VPWR VGND sg13g2_decap_8
XFILLER_33_614 VPWR VGND sg13g2_decap_8
XFILLER_14_850 VPWR VGND sg13g2_decap_8
XFILLER_32_124 VPWR VGND sg13g2_decap_8
XFILLER_20_319 VPWR VGND sg13g2_decap_8
XFILLER_41_691 VPWR VGND sg13g2_decap_8
XFILLER_13_382 VPWR VGND sg13g2_decap_8
XFILLER_9_375 VPWR VGND sg13g2_decap_8
XFILLER_5_592 VPWR VGND sg13g2_decap_8
XFILLER_49_791 VPWR VGND sg13g2_decap_8
XFILLER_36_452 VPWR VGND sg13g2_decap_8
XFILLER_37_986 VPWR VGND sg13g2_decap_8
XFILLER_23_102 VPWR VGND sg13g2_decap_8
XFILLER_12_809 VPWR VGND sg13g2_decap_8
XFILLER_24_669 VPWR VGND sg13g2_decap_8
XFILLER_11_319 VPWR VGND sg13g2_decap_8
XFILLER_20_831 VPWR VGND sg13g2_decap_8
XFILLER_32_691 VPWR VGND sg13g2_decap_8
XFILLER_11_46 VPWR VGND sg13g2_decap_8
XFILLER_3_529 VPWR VGND sg13g2_decap_8
XFILLER_47_728 VPWR VGND sg13g2_decap_8
XFILLER_19_419 VPWR VGND sg13g2_decap_8
XFILLER_46_238 VPWR VGND sg13g2_decap_8
XFILLER_28_953 VPWR VGND sg13g2_decap_8
XFILLER_43_901 VPWR VGND sg13g2_decap_8
XFILLER_27_441 VPWR VGND sg13g2_decap_8
XFILLER_36_54 VPWR VGND sg13g2_decap_8
XFILLER_39_290 VPWR VGND sg13g2_decap_8
XFILLER_42_411 VPWR VGND sg13g2_decap_8
XFILLER_14_102 VPWR VGND sg13g2_decap_8
XFILLER_43_978 VPWR VGND sg13g2_decap_8
XFILLER_15_658 VPWR VGND sg13g2_decap_8
XFILLER_42_488 VPWR VGND sg13g2_decap_8
XFILLER_14_179 VPWR VGND sg13g2_decap_8
XFILLER_35_1011 VPWR VGND sg13g2_decap_8
XFILLER_30_639 VPWR VGND sg13g2_decap_8
XFILLER_11_886 VPWR VGND sg13g2_decap_8
XFILLER_7_868 VPWR VGND sg13g2_decap_8
XFILLER_6_312 VPWR VGND sg13g2_decap_8
XFILLER_10_396 VPWR VGND sg13g2_decap_8
XFILLER_6_389 VPWR VGND sg13g2_decap_8
XFILLER_18_452 VPWR VGND sg13g2_decap_8
XFILLER_19_986 VPWR VGND sg13g2_decap_8
XFILLER_45_271 VPWR VGND sg13g2_decap_8
XFILLER_34_923 VPWR VGND sg13g2_decap_8
XFILLER_33_488 VPWR VGND sg13g2_decap_8
XFILLER_20_116 VPWR VGND sg13g2_decap_8
XFILLER_9_172 VPWR VGND sg13g2_decap_8
XFILLER_29_739 VPWR VGND sg13g2_decap_8
XFILLER_25_901 VPWR VGND sg13g2_decap_8
XFILLER_43_208 VPWR VGND sg13g2_decap_8
XFILLER_37_783 VPWR VGND sg13g2_decap_8
XFILLER_25_978 VPWR VGND sg13g2_decap_8
XFILLER_36_282 VPWR VGND sg13g2_decap_4
XFILLER_12_606 VPWR VGND sg13g2_decap_8
XFILLER_19_1028 VPWR VGND sg13g2_fill_1
XFILLER_24_466 VPWR VGND sg13g2_decap_8
XFILLER_40_915 VPWR VGND sg13g2_decap_8
XFILLER_11_116 VPWR VGND sg13g2_decap_8
XFILLER_22_67 VPWR VGND sg13g2_decap_8
XFILLER_4_816 VPWR VGND sg13g2_decap_8
XFILLER_3_326 VPWR VGND sg13g2_decap_8
XFILLER_47_525 VPWR VGND sg13g2_decap_8
XFILLER_47_42 VPWR VGND sg13g2_decap_8
XFILLER_19_227 VPWR VGND sg13g2_decap_8
XFILLER_28_750 VPWR VGND sg13g2_decap_8
XFILLER_16_923 VPWR VGND sg13g2_decap_8
XFILLER_43_775 VPWR VGND sg13g2_decap_8
XFILLER_15_455 VPWR VGND sg13g2_decap_8
XFILLER_31_904 VPWR VGND sg13g2_decap_8
XFILLER_42_285 VPWR VGND sg13g2_decap_8
XFILLER_30_436 VPWR VGND sg13g2_decap_8
XFILLER_8_25 VPWR VGND sg13g2_decap_8
XFILLER_11_683 VPWR VGND sg13g2_decap_8
XFILLER_10_193 VPWR VGND sg13g2_decap_8
XFILLER_7_665 VPWR VGND sg13g2_decap_8
X_157_ net29 net25 VPWR VGND sg13g2_buf_1
XFILLER_6_186 VPWR VGND sg13g2_decap_8
X_088_ _053_ mod1.i_out_qam16\[3\] net11 VPWR VGND sg13g2_nand2_1
XFILLER_3_893 VPWR VGND sg13g2_decap_8
XFILLER_33_5 VPWR VGND sg13g2_decap_8
XFILLER_26_4 VPWR VGND sg13g2_decap_8
XFILLER_38_547 VPWR VGND sg13g2_decap_8
XFILLER_19_783 VPWR VGND sg13g2_decap_8
XFILLER_34_720 VPWR VGND sg13g2_decap_8
XFILLER_22_926 VPWR VGND sg13g2_decap_8
XFILLER_34_797 VPWR VGND sg13g2_decap_8
XFILLER_21_458 VPWR VGND sg13g2_decap_8
XFILLER_1_819 VPWR VGND sg13g2_decap_8
XFILLER_0_329 VPWR VGND sg13g2_decap_8
XFILLER_29_536 VPWR VGND sg13g2_decap_8
XFILLER_17_56 VPWR VGND sg13g2_decap_8
XFILLER_37_580 VPWR VGND sg13g2_decap_8
XFILLER_12_403 VPWR VGND sg13g2_decap_8
XFILLER_25_775 VPWR VGND sg13g2_decap_8
XFILLER_40_712 VPWR VGND sg13g2_decap_8
XFILLER_24_285 VPWR VGND sg13g2_decap_8
XFILLER_33_33 VPWR VGND sg13g2_decap_8
XFILLER_40_789 VPWR VGND sg13g2_decap_8
XFILLER_4_613 VPWR VGND sg13g2_decap_8
XFILLER_3_123 VPWR VGND sg13g2_decap_8
XFILLER_48_812 VPWR VGND sg13g2_decap_8
XFILLER_47_322 VPWR VGND sg13g2_decap_8
XFILLER_0_896 VPWR VGND sg13g2_decap_8
XFILLER_48_889 VPWR VGND sg13g2_decap_8
XFILLER_35_528 VPWR VGND sg13g2_decap_8
XFILLER_47_399 VPWR VGND sg13g2_decap_8
XFILLER_16_720 VPWR VGND sg13g2_decap_8
XFILLER_31_701 VPWR VGND sg13g2_decap_8
XFILLER_43_572 VPWR VGND sg13g2_decap_8
XFILLER_16_797 VPWR VGND sg13g2_decap_8
XFILLER_30_222 VPWR VGND sg13g2_decap_8
XFILLER_31_778 VPWR VGND sg13g2_decap_8
XFILLER_12_970 VPWR VGND sg13g2_decap_8
XFILLER_8_963 VPWR VGND sg13g2_decap_8
XFILLER_11_480 VPWR VGND sg13g2_decap_8
XFILLER_7_462 VPWR VGND sg13g2_decap_8
XFILLER_3_690 VPWR VGND sg13g2_decap_8
XFILLER_39_823 VPWR VGND sg13g2_decap_8
XFILLER_17_0 VPWR VGND sg13g2_decap_8
XFILLER_38_333 VPWR VGND sg13g2_decap_8
XFILLER_0_1001 VPWR VGND sg13g2_decap_8
XFILLER_0_70 VPWR VGND sg13g2_decap_8
XFILLER_19_580 VPWR VGND sg13g2_decap_8
XFILLER_26_539 VPWR VGND sg13g2_decap_8
XFILLER_41_509 VPWR VGND sg13g2_decap_8
XFILLER_21_211 VPWR VGND sg13g2_decap_8
XFILLER_22_723 VPWR VGND sg13g2_decap_8
XFILLER_34_594 VPWR VGND sg13g2_decap_8
XFILLER_10_907 VPWR VGND sg13g2_decap_8
XFILLER_21_222 VPWR VGND sg13g2_fill_1
XFILLER_21_277 VPWR VGND sg13g2_decap_8
XFILLER_1_616 VPWR VGND sg13g2_decap_8
XFILLER_0_126 VPWR VGND sg13g2_decap_8
XFILLER_49_609 VPWR VGND sg13g2_decap_8
XFILLER_48_119 VPWR VGND sg13g2_decap_8
XFILLER_28_11 VPWR VGND sg13g2_decap_8
XFILLER_28_88 VPWR VGND sg13g2_decap_8
XFILLER_45_859 VPWR VGND sg13g2_decap_8
XFILLER_17_539 VPWR VGND sg13g2_decap_8
XFILLER_44_369 VPWR VGND sg13g2_decap_8
XFILLER_32_509 VPWR VGND sg13g2_decap_8
XFILLER_44_54 VPWR VGND sg13g2_decap_8
XFILLER_12_200 VPWR VGND sg13g2_decap_8
XFILLER_25_572 VPWR VGND sg13g2_decap_8
XFILLER_13_767 VPWR VGND sg13g2_decap_8
XFILLER_12_277 VPWR VGND sg13g2_decap_8
XFILLER_40_586 VPWR VGND sg13g2_decap_8
XFILLER_5_900 VPWR VGND sg13g2_decap_8
XFILLER_4_410 VPWR VGND sg13g2_decap_8
XFILLER_5_977 VPWR VGND sg13g2_decap_8
XFILLER_4_487 VPWR VGND sg13g2_decap_8
XFILLER_0_693 VPWR VGND sg13g2_decap_8
XFILLER_48_686 VPWR VGND sg13g2_decap_8
XFILLER_36_837 VPWR VGND sg13g2_decap_8
XFILLER_47_196 VPWR VGND sg13g2_decap_8
XFILLER_35_325 VPWR VGND sg13g2_decap_8
XFILLER_16_594 VPWR VGND sg13g2_decap_8
XFILLER_31_575 VPWR VGND sg13g2_decap_8
XFILLER_8_760 VPWR VGND sg13g2_decap_8
XFILLER_39_620 VPWR VGND sg13g2_decap_8
XFILLER_22_1024 VPWR VGND sg13g2_decap_4
XFILLER_38_130 VPWR VGND sg13g2_decap_8
XFILLER_27_826 VPWR VGND sg13g2_decap_8
XFILLER_26_336 VPWR VGND sg13g2_decap_8
XFILLER_39_697 VPWR VGND sg13g2_decap_8
XFILLER_41_306 VPWR VGND sg13g2_decap_8
XFILLER_22_520 VPWR VGND sg13g2_decap_8
XFILLER_35_892 VPWR VGND sg13g2_decap_8
XFILLER_34_391 VPWR VGND sg13g2_decap_8
XFILLER_10_704 VPWR VGND sg13g2_decap_8
XFILLER_14_46 VPWR VGND sg13g2_decap_8
XFILLER_22_597 VPWR VGND sg13g2_decap_8
XFILLER_5_207 VPWR VGND sg13g2_decap_8
XFILLER_30_12 VPWR VGND sg13g2_decap_8
XFILLER_2_914 VPWR VGND sg13g2_decap_8
XFILLER_30_89 VPWR VGND sg13g2_decap_8
XFILLER_1_413 VPWR VGND sg13g2_decap_8
XFILLER_49_406 VPWR VGND sg13g2_decap_8
XFILLER_39_32 VPWR VGND sg13g2_decap_8
XFILLER_17_336 VPWR VGND sg13g2_decap_8
XFILLER_18_837 VPWR VGND sg13g2_decap_8
XFILLER_45_656 VPWR VGND sg13g2_decap_8
XFILLER_44_166 VPWR VGND sg13g2_decap_8
XFILLER_32_306 VPWR VGND sg13g2_decap_8
XFILLER_41_873 VPWR VGND sg13g2_decap_8
XFILLER_13_564 VPWR VGND sg13g2_decap_8
XFILLER_9_557 VPWR VGND sg13g2_decap_8
XFILLER_40_383 VPWR VGND sg13g2_decap_8
XFILLER_5_774 VPWR VGND sg13g2_decap_8
XFILLER_4_284 VPWR VGND sg13g2_decap_8
XFILLER_45_1013 VPWR VGND sg13g2_decap_8
XFILLER_1_980 VPWR VGND sg13g2_decap_8
XFILLER_0_490 VPWR VGND sg13g2_decap_8
XFILLER_49_973 VPWR VGND sg13g2_decap_8
XFILLER_48_483 VPWR VGND sg13g2_decap_8
XFILLER_36_634 VPWR VGND sg13g2_decap_8
XFILLER_35_166 VPWR VGND sg13g2_decap_8
XFILLER_16_391 VPWR VGND sg13g2_decap_8
XFILLER_35_199 VPWR VGND sg13g2_fill_2
XFILLER_32_873 VPWR VGND sg13g2_decap_8
XFILLER_31_372 VPWR VGND sg13g2_decap_8
XFILLER_27_623 VPWR VGND sg13g2_decap_8
XFILLER_39_494 VPWR VGND sg13g2_decap_8
XFILLER_26_144 VPWR VGND sg13g2_decap_8
XFILLER_14_339 VPWR VGND sg13g2_decap_8
XFILLER_23_851 VPWR VGND sg13g2_decap_8
XFILLER_25_67 VPWR VGND sg13g2_decap_8
XFILLER_10_501 VPWR VGND sg13g2_decap_8
XFILLER_41_158 VPWR VGND sg13g2_decap_8
XFILLER_22_383 VPWR VGND sg13g2_decap_4
XFILLER_41_11 VPWR VGND sg13g2_decap_8
XFILLER_10_578 VPWR VGND sg13g2_decap_8
XFILLER_41_88 VPWR VGND sg13g2_decap_8
XFILLER_2_711 VPWR VGND sg13g2_decap_8
XFILLER_1_210 VPWR VGND sg13g2_decap_8
XFILLER_29_1019 VPWR VGND sg13g2_decap_8
XFILLER_49_203 VPWR VGND sg13g2_decap_8
XFILLER_2_788 VPWR VGND sg13g2_decap_8
XFILLER_1_287 VPWR VGND sg13g2_decap_8
XFILLER_46_910 VPWR VGND sg13g2_decap_8
XFILLER_18_634 VPWR VGND sg13g2_decap_8
XFILLER_46_987 VPWR VGND sg13g2_decap_8
XFILLER_45_453 VPWR VGND sg13g2_decap_8
XFILLER_17_133 VPWR VGND sg13g2_decap_8
XFILLER_32_103 VPWR VGND sg13g2_decap_8
XFILLER_41_670 VPWR VGND sg13g2_decap_8
XFILLER_13_361 VPWR VGND sg13g2_decap_8
XFILLER_9_354 VPWR VGND sg13g2_decap_8
XFILLER_12_1012 VPWR VGND sg13g2_decap_8
XFILLER_5_571 VPWR VGND sg13g2_decap_8
XFILLER_49_770 VPWR VGND sg13g2_decap_8
XFILLER_48_280 VPWR VGND sg13g2_decap_8
XFILLER_36_431 VPWR VGND sg13g2_decap_8
XFILLER_37_965 VPWR VGND sg13g2_decap_8
XFILLER_24_648 VPWR VGND sg13g2_decap_8
XFILLER_20_810 VPWR VGND sg13g2_decap_8
XFILLER_23_158 VPWR VGND sg13g2_decap_8
XFILLER_32_670 VPWR VGND sg13g2_decap_8
XFILLER_31_180 VPWR VGND sg13g2_decap_8
XFILLER_20_887 VPWR VGND sg13g2_decap_8
XFILLER_3_508 VPWR VGND sg13g2_decap_8
XFILLER_11_25 VPWR VGND sg13g2_decap_8
XFILLER_47_707 VPWR VGND sg13g2_decap_8
XFILLER_46_217 VPWR VGND sg13g2_decap_8
XFILLER_27_420 VPWR VGND sg13g2_decap_8
XFILLER_28_932 VPWR VGND sg13g2_decap_8
XFILLER_36_33 VPWR VGND sg13g2_decap_8
XFILLER_43_957 VPWR VGND sg13g2_decap_8
XFILLER_15_637 VPWR VGND sg13g2_decap_8
XFILLER_27_497 VPWR VGND sg13g2_decap_8
XFILLER_42_467 VPWR VGND sg13g2_decap_8
XFILLER_14_158 VPWR VGND sg13g2_decap_8
XFILLER_30_618 VPWR VGND sg13g2_decap_8
XFILLER_11_865 VPWR VGND sg13g2_decap_8
XFILLER_22_180 VPWR VGND sg13g2_decap_8
XFILLER_10_375 VPWR VGND sg13g2_decap_8
XFILLER_7_847 VPWR VGND sg13g2_decap_8
XFILLER_6_368 VPWR VGND sg13g2_decap_8
XFILLER_2_585 VPWR VGND sg13g2_decap_8
XFILLER_42_1027 VPWR VGND sg13g2_fill_2
XFILLER_38_729 VPWR VGND sg13g2_decap_8
XFILLER_18_431 VPWR VGND sg13g2_decap_8
XFILLER_19_965 VPWR VGND sg13g2_decap_8
XFILLER_34_902 VPWR VGND sg13g2_decap_8
XFILLER_46_784 VPWR VGND sg13g2_decap_8
XFILLER_45_250 VPWR VGND sg13g2_decap_8
XFILLER_34_979 VPWR VGND sg13g2_decap_8
XFILLER_33_467 VPWR VGND sg13g2_decap_8
XFILLER_9_151 VPWR VGND sg13g2_decap_8
XFILLER_47_0 VPWR VGND sg13g2_decap_8
XFILLER_3_81 VPWR VGND sg13g2_decap_8
XFILLER_29_718 VPWR VGND sg13g2_decap_8
XFILLER_28_239 VPWR VGND sg13g2_decap_4
XFILLER_36_261 VPWR VGND sg13g2_decap_8
XFILLER_37_762 VPWR VGND sg13g2_decap_8
XFILLER_19_1007 VPWR VGND sg13g2_decap_8
XFILLER_24_445 VPWR VGND sg13g2_decap_8
XFILLER_25_957 VPWR VGND sg13g2_decap_8
XFILLER_20_684 VPWR VGND sg13g2_decap_8
XFILLER_22_46 VPWR VGND sg13g2_decap_8
XFILLER_3_305 VPWR VGND sg13g2_decap_8
XFILLER_47_504 VPWR VGND sg13g2_decap_8
XFILLER_47_21 VPWR VGND sg13g2_decap_8
XFILLER_19_206 VPWR VGND sg13g2_decap_8
XFILLER_47_98 VPWR VGND sg13g2_decap_8
XFILLER_16_902 VPWR VGND sg13g2_decap_8
XFILLER_43_754 VPWR VGND sg13g2_decap_8
XFILLER_15_434 VPWR VGND sg13g2_decap_8
XFILLER_42_264 VPWR VGND sg13g2_decap_8
XFILLER_16_979 VPWR VGND sg13g2_decap_8
XFILLER_30_415 VPWR VGND sg13g2_decap_8
XFILLER_11_662 VPWR VGND sg13g2_decap_8
XFILLER_10_172 VPWR VGND sg13g2_decap_8
XFILLER_7_644 VPWR VGND sg13g2_decap_8
XFILLER_6_165 VPWR VGND sg13g2_decap_8
X_087_ _050_ _051_ _049_ net27 VPWR VGND _052_ sg13g2_nand4_1
XFILLER_3_872 VPWR VGND sg13g2_decap_8
XFILLER_2_382 VPWR VGND sg13g2_decap_8
XFILLER_19_4 VPWR VGND sg13g2_decap_8
XFILLER_38_526 VPWR VGND sg13g2_decap_8
XFILLER_19_762 VPWR VGND sg13g2_decap_8
XFILLER_46_581 VPWR VGND sg13g2_decap_8
XFILLER_22_905 VPWR VGND sg13g2_decap_8
XFILLER_34_776 VPWR VGND sg13g2_decap_8
XFILLER_21_437 VPWR VGND sg13g2_decap_8
XFILLER_30_982 VPWR VGND sg13g2_decap_8
XFILLER_0_308 VPWR VGND sg13g2_decap_8
XFILLER_29_515 VPWR VGND sg13g2_decap_8
XFILLER_17_35 VPWR VGND sg13g2_decap_8
XFILLER_25_754 VPWR VGND sg13g2_decap_8
XFILLER_13_949 VPWR VGND sg13g2_decap_8
XFILLER_24_264 VPWR VGND sg13g2_decap_8
XFILLER_33_12 VPWR VGND sg13g2_decap_8
XFILLER_12_459 VPWR VGND sg13g2_decap_8
XFILLER_40_768 VPWR VGND sg13g2_decap_8
XFILLER_33_89 VPWR VGND sg13g2_decap_8
XFILLER_20_481 VPWR VGND sg13g2_decap_8
XFILLER_3_102 VPWR VGND sg13g2_decap_8
XFILLER_4_669 VPWR VGND sg13g2_decap_8
XFILLER_3_179 VPWR VGND sg13g2_decap_8
XFILLER_0_875 VPWR VGND sg13g2_decap_8
XFILLER_47_301 VPWR VGND sg13g2_decap_8
XFILLER_48_868 VPWR VGND sg13g2_decap_8
XFILLER_47_378 VPWR VGND sg13g2_decap_8
XFILLER_35_507 VPWR VGND sg13g2_decap_8
XFILLER_43_551 VPWR VGND sg13g2_decap_8
XFILLER_16_776 VPWR VGND sg13g2_decap_8
XFILLER_30_201 VPWR VGND sg13g2_decap_8
XFILLER_31_757 VPWR VGND sg13g2_decap_8
XFILLER_30_278 VPWR VGND sg13g2_decap_8
XFILLER_8_942 VPWR VGND sg13g2_decap_8
XFILLER_7_441 VPWR VGND sg13g2_decap_8
X_139_ net15 VGND VPWR _002_ Demo1.epsk_de1.bit_out\[1\] clknet_2_3__leaf_clk sg13g2_dfrbpq_1
XFILLER_48_1022 VPWR VGND sg13g2_decap_8
XFILLER_39_802 VPWR VGND sg13g2_decap_8
XFILLER_38_312 VPWR VGND sg13g2_decap_8
XFILLER_39_879 VPWR VGND sg13g2_decap_8
XFILLER_26_518 VPWR VGND sg13g2_decap_8
XFILLER_22_702 VPWR VGND sg13g2_decap_8
XFILLER_34_573 VPWR VGND sg13g2_decap_8
XFILLER_21_256 VPWR VGND sg13g2_decap_8
XFILLER_22_779 VPWR VGND sg13g2_decap_8
XFILLER_0_105 VPWR VGND sg13g2_decap_8
XFILLER_29_345 VPWR VGND sg13g2_fill_2
XFILLER_45_838 VPWR VGND sg13g2_decap_8
XFILLER_17_518 VPWR VGND sg13g2_decap_8
XFILLER_28_67 VPWR VGND sg13g2_decap_8
XFILLER_44_348 VPWR VGND sg13g2_decap_8
XFILLER_29_389 VPWR VGND sg13g2_decap_8
XFILLER_38_890 VPWR VGND sg13g2_decap_8
XFILLER_44_33 VPWR VGND sg13g2_decap_8
XFILLER_25_551 VPWR VGND sg13g2_decap_8
XFILLER_13_746 VPWR VGND sg13g2_decap_8
XFILLER_9_739 VPWR VGND sg13g2_decap_8
XFILLER_12_256 VPWR VGND sg13g2_decap_8
XFILLER_40_565 VPWR VGND sg13g2_decap_8
XFILLER_8_249 VPWR VGND sg13g2_decap_8
XFILLER_5_956 VPWR VGND sg13g2_decap_8
XFILLER_4_466 VPWR VGND sg13g2_decap_8
XFILLER_0_672 VPWR VGND sg13g2_decap_8
XFILLER_39_109 VPWR VGND sg13g2_decap_8
XFILLER_48_665 VPWR VGND sg13g2_decap_8
Xclkbuf_2_3__f_clk clknet_0_clk clknet_2_3__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_35_304 VPWR VGND sg13g2_decap_8
XFILLER_36_816 VPWR VGND sg13g2_decap_8
XFILLER_47_175 VPWR VGND sg13g2_decap_8
XFILLER_16_573 VPWR VGND sg13g2_decap_8
XFILLER_31_554 VPWR VGND sg13g2_decap_8
XFILLER_22_1003 VPWR VGND sg13g2_decap_8
XFILLER_26_304 VPWR VGND sg13g2_decap_4
XFILLER_27_805 VPWR VGND sg13g2_decap_8
XFILLER_39_676 VPWR VGND sg13g2_decap_8
XFILLER_38_186 VPWR VGND sg13g2_decap_8
XFILLER_35_871 VPWR VGND sg13g2_decap_8
XFILLER_14_25 VPWR VGND sg13g2_decap_8
XFILLER_22_576 VPWR VGND sg13g2_decap_8
XFILLER_30_68 VPWR VGND sg13g2_decap_8
XFILLER_7_1008 VPWR VGND sg13g2_decap_8
XFILLER_39_11 VPWR VGND sg13g2_decap_8
XFILLER_1_469 VPWR VGND sg13g2_decap_8
XFILLER_39_88 VPWR VGND sg13g2_decap_8
XFILLER_18_816 VPWR VGND sg13g2_decap_8
XFILLER_45_635 VPWR VGND sg13g2_decap_8
XFILLER_17_315 VPWR VGND sg13g2_decap_8
XFILLER_29_175 VPWR VGND sg13g2_decap_8
XFILLER_44_145 VPWR VGND sg13g2_decap_8
XFILLER_26_882 VPWR VGND sg13g2_decap_8
XFILLER_41_852 VPWR VGND sg13g2_decap_8
XFILLER_13_543 VPWR VGND sg13g2_decap_8
XFILLER_25_381 VPWR VGND sg13g2_decap_8
XFILLER_40_362 VPWR VGND sg13g2_decap_8
XFILLER_9_536 VPWR VGND sg13g2_decap_8
XFILLER_5_753 VPWR VGND sg13g2_decap_8
XFILLER_4_263 VPWR VGND sg13g2_decap_8
XFILLER_49_952 VPWR VGND sg13g2_decap_8
XFILLER_48_462 VPWR VGND sg13g2_decap_8
XFILLER_36_613 VPWR VGND sg13g2_decap_8
XFILLER_35_145 VPWR VGND sg13g2_decap_8
XFILLER_17_882 VPWR VGND sg13g2_decap_8
XFILLER_16_370 VPWR VGND sg13g2_decap_8
XFILLER_32_852 VPWR VGND sg13g2_decap_8
XFILLER_31_351 VPWR VGND sg13g2_decap_8
XFILLER_6_81 VPWR VGND sg13g2_decap_8
XFILLER_27_602 VPWR VGND sg13g2_decap_8
XFILLER_39_473 VPWR VGND sg13g2_decap_8
XFILLER_15_819 VPWR VGND sg13g2_decap_8
XFILLER_26_123 VPWR VGND sg13g2_decap_8
XFILLER_27_679 VPWR VGND sg13g2_decap_8
XFILLER_14_318 VPWR VGND sg13g2_decap_8
XFILLER_42_649 VPWR VGND sg13g2_decap_8
XFILLER_23_830 VPWR VGND sg13g2_decap_8
XFILLER_25_46 VPWR VGND sg13g2_decap_8
XFILLER_41_137 VPWR VGND sg13g2_decap_8
XFILLER_22_362 VPWR VGND sg13g2_decap_8
XFILLER_10_557 VPWR VGND sg13g2_decap_8
XFILLER_41_67 VPWR VGND sg13g2_decap_8
XFILLER_2_767 VPWR VGND sg13g2_decap_8
XFILLER_1_266 VPWR VGND sg13g2_decap_8
XFILLER_2_39 VPWR VGND sg13g2_decap_8
XFILLER_49_259 VPWR VGND sg13g2_decap_8
XFILLER_17_112 VPWR VGND sg13g2_decap_8
XFILLER_18_613 VPWR VGND sg13g2_decap_8
XFILLER_46_966 VPWR VGND sg13g2_decap_8
XFILLER_45_432 VPWR VGND sg13g2_decap_8
XFILLER_17_189 VPWR VGND sg13g2_decap_8
XFILLER_33_649 VPWR VGND sg13g2_decap_8
XFILLER_13_340 VPWR VGND sg13g2_decap_8
XFILLER_14_885 VPWR VGND sg13g2_decap_8
XFILLER_32_159 VPWR VGND sg13g2_decap_8
XFILLER_9_333 VPWR VGND sg13g2_decap_8
XFILLER_5_550 VPWR VGND sg13g2_decap_8
XFILLER_36_410 VPWR VGND sg13g2_decap_8
XFILLER_37_944 VPWR VGND sg13g2_decap_8
XFILLER_24_627 VPWR VGND sg13g2_decap_8
XFILLER_36_487 VPWR VGND sg13g2_decap_8
XFILLER_23_137 VPWR VGND sg13g2_decap_8
XFILLER_20_866 VPWR VGND sg13g2_decap_8
XFILLER_28_911 VPWR VGND sg13g2_decap_8
XFILLER_36_12 VPWR VGND sg13g2_decap_8
XFILLER_39_270 VPWR VGND sg13g2_decap_8
XFILLER_43_936 VPWR VGND sg13g2_decap_8
XFILLER_15_616 VPWR VGND sg13g2_decap_8
XFILLER_27_476 VPWR VGND sg13g2_decap_8
XFILLER_28_988 VPWR VGND sg13g2_decap_8
XFILLER_42_446 VPWR VGND sg13g2_decap_8
XFILLER_14_137 VPWR VGND sg13g2_decap_8
XFILLER_36_89 VPWR VGND sg13g2_decap_8
XFILLER_11_844 VPWR VGND sg13g2_decap_8
XFILLER_10_354 VPWR VGND sg13g2_decap_8
XFILLER_7_826 VPWR VGND sg13g2_decap_8
XFILLER_6_347 VPWR VGND sg13g2_decap_8
XFILLER_7_0 VPWR VGND sg13g2_decap_8
XFILLER_2_564 VPWR VGND sg13g2_decap_8
XFILLER_42_1006 VPWR VGND sg13g2_decap_8
XFILLER_38_708 VPWR VGND sg13g2_decap_8
XFILLER_18_410 VPWR VGND sg13g2_decap_8
XFILLER_37_229 VPWR VGND sg13g2_decap_8
XFILLER_19_944 VPWR VGND sg13g2_decap_8
XFILLER_46_763 VPWR VGND sg13g2_decap_8
XFILLER_18_487 VPWR VGND sg13g2_decap_8
XFILLER_33_446 VPWR VGND sg13g2_decap_8
XFILLER_34_958 VPWR VGND sg13g2_decap_8
XFILLER_21_619 VPWR VGND sg13g2_decap_8
XFILLER_14_682 VPWR VGND sg13g2_decap_8
XFILLER_9_130 VPWR VGND sg13g2_decap_8
XFILLER_3_60 VPWR VGND sg13g2_decap_8
XFILLER_28_218 VPWR VGND sg13g2_decap_8
XFILLER_37_741 VPWR VGND sg13g2_decap_8
XFILLER_36_240 VPWR VGND sg13g2_decap_8
XFILLER_24_424 VPWR VGND sg13g2_decap_8
XFILLER_25_936 VPWR VGND sg13g2_decap_8
XFILLER_22_25 VPWR VGND sg13g2_decap_8
XFILLER_20_663 VPWR VGND sg13g2_decap_8
XFILLER_0_7 VPWR VGND sg13g2_decap_8
XFILLER_47_77 VPWR VGND sg13g2_decap_8
XFILLER_28_785 VPWR VGND sg13g2_decap_8
XFILLER_43_733 VPWR VGND sg13g2_decap_8
XFILLER_15_413 VPWR VGND sg13g2_decap_8
XFILLER_16_958 VPWR VGND sg13g2_decap_8
XFILLER_27_273 VPWR VGND sg13g2_decap_8
XFILLER_42_243 VPWR VGND sg13g2_decap_8
XFILLER_24_991 VPWR VGND sg13g2_decap_8
XFILLER_31_939 VPWR VGND sg13g2_decap_8
XFILLER_11_641 VPWR VGND sg13g2_decap_8
XFILLER_10_151 VPWR VGND sg13g2_decap_8
XFILLER_7_623 VPWR VGND sg13g2_decap_8
XFILLER_6_144 VPWR VGND sg13g2_decap_8
X_086_ _052_ mod1.i_out_qam16\[2\] net11 VPWR VGND sg13g2_nand2_1
XFILLER_3_851 VPWR VGND sg13g2_decap_8
XFILLER_2_361 VPWR VGND sg13g2_decap_8
XFILLER_38_505 VPWR VGND sg13g2_decap_8
XFILLER_19_741 VPWR VGND sg13g2_decap_8
XFILLER_46_560 VPWR VGND sg13g2_decap_8
XFILLER_18_284 VPWR VGND sg13g2_decap_8
XFILLER_33_210 VPWR VGND sg13g2_decap_8
XFILLER_33_243 VPWR VGND sg13g2_decap_8
XFILLER_34_755 VPWR VGND sg13g2_decap_8
XFILLER_15_980 VPWR VGND sg13g2_decap_8
XFILLER_21_416 VPWR VGND sg13g2_decap_8
XFILLER_33_298 VPWR VGND sg13g2_decap_8
XFILLER_30_961 VPWR VGND sg13g2_decap_8
XFILLER_17_14 VPWR VGND sg13g2_decap_8
XFILLER_25_733 VPWR VGND sg13g2_decap_8
XFILLER_24_243 VPWR VGND sg13g2_decap_8
XFILLER_13_928 VPWR VGND sg13g2_decap_8
XFILLER_12_438 VPWR VGND sg13g2_decap_8
XFILLER_33_68 VPWR VGND sg13g2_decap_8
XFILLER_40_747 VPWR VGND sg13g2_decap_8
XFILLER_20_460 VPWR VGND sg13g2_decap_8
XFILLER_21_983 VPWR VGND sg13g2_decap_8
XFILLER_32_1027 VPWR VGND sg13g2_fill_2
XFILLER_4_648 VPWR VGND sg13g2_decap_8
XFILLER_3_158 VPWR VGND sg13g2_decap_8
XFILLER_0_854 VPWR VGND sg13g2_decap_8
XFILLER_48_847 VPWR VGND sg13g2_decap_8
XFILLER_47_357 VPWR VGND sg13g2_decap_8
XFILLER_28_582 VPWR VGND sg13g2_decap_8
XFILLER_43_530 VPWR VGND sg13g2_decap_8
XFILLER_16_755 VPWR VGND sg13g2_decap_8
XFILLER_15_254 VPWR VGND sg13g2_decap_8
XFILLER_31_736 VPWR VGND sg13g2_decap_8
XFILLER_8_921 VPWR VGND sg13g2_decap_8
XFILLER_30_257 VPWR VGND sg13g2_decap_8
XFILLER_7_420 VPWR VGND sg13g2_decap_8
XFILLER_8_998 VPWR VGND sg13g2_decap_8
X_138_ net14 VGND VPWR _001_ Demo1.epsk_de1.bit_out\[0\] clknet_2_1__leaf_clk sg13g2_dfrbpq_1
XFILLER_48_1001 VPWR VGND sg13g2_decap_8
XFILLER_7_497 VPWR VGND sg13g2_decap_8
X_069_ _042_ _041_ Demo1.epsk_de1.bit_out\[0\] net11 Demo1.qam16_bits\[0\] VPWR VGND
+ sg13g2_a22oi_1
XFILLER_39_858 VPWR VGND sg13g2_decap_8
XFILLER_38_368 VPWR VGND sg13g2_decap_4
XFILLER_38_379 VPWR VGND sg13g2_decap_8
XFILLER_34_552 VPWR VGND sg13g2_decap_8
XFILLER_21_235 VPWR VGND sg13g2_decap_8
XFILLER_22_758 VPWR VGND sg13g2_decap_8
XFILLER_9_81 VPWR VGND sg13g2_decap_8
XFILLER_28_46 VPWR VGND sg13g2_decap_8
XFILLER_29_324 VPWR VGND sg13g2_decap_8
XFILLER_45_817 VPWR VGND sg13g2_decap_8
XFILLER_44_327 VPWR VGND sg13g2_decap_8
XFILLER_44_12 VPWR VGND sg13g2_decap_8
XFILLER_25_530 VPWR VGND sg13g2_decap_8
XFILLER_13_725 VPWR VGND sg13g2_decap_8
XFILLER_44_89 VPWR VGND sg13g2_decap_8
XFILLER_9_718 VPWR VGND sg13g2_decap_8
XFILLER_12_235 VPWR VGND sg13g2_decap_8
XFILLER_40_544 VPWR VGND sg13g2_decap_8
XFILLER_8_228 VPWR VGND sg13g2_decap_8
XFILLER_21_780 VPWR VGND sg13g2_decap_8
XFILLER_5_935 VPWR VGND sg13g2_decap_8
XFILLER_5_39 VPWR VGND sg13g2_decap_8
XFILLER_4_445 VPWR VGND sg13g2_decap_8
XFILLER_0_651 VPWR VGND sg13g2_decap_8
XFILLER_48_644 VPWR VGND sg13g2_decap_8
XFILLER_47_154 VPWR VGND sg13g2_decap_8
XFILLER_16_552 VPWR VGND sg13g2_decap_8
XFILLER_44_894 VPWR VGND sg13g2_decap_8
XFILLER_31_533 VPWR VGND sg13g2_decap_8
XFILLER_15_1022 VPWR VGND sg13g2_decap_8
XFILLER_8_795 VPWR VGND sg13g2_decap_8
XFILLER_7_294 VPWR VGND sg13g2_decap_8
XFILLER_39_655 VPWR VGND sg13g2_decap_8
XFILLER_38_165 VPWR VGND sg13g2_decap_8
XFILLER_35_850 VPWR VGND sg13g2_decap_8
XFILLER_22_555 VPWR VGND sg13g2_decap_8
XFILLER_10_739 VPWR VGND sg13g2_decap_8
XFILLER_30_47 VPWR VGND sg13g2_decap_8
XFILLER_2_949 VPWR VGND sg13g2_decap_8
XFILLER_1_448 VPWR VGND sg13g2_decap_8
XFILLER_39_67 VPWR VGND sg13g2_decap_8
XFILLER_29_154 VPWR VGND sg13g2_decap_8
XFILLER_45_614 VPWR VGND sg13g2_decap_8
XFILLER_44_124 VPWR VGND sg13g2_decap_8
XFILLER_25_360 VPWR VGND sg13g2_decap_8
XFILLER_26_861 VPWR VGND sg13g2_decap_8
XFILLER_41_831 VPWR VGND sg13g2_decap_8
XFILLER_13_522 VPWR VGND sg13g2_decap_8
XFILLER_9_515 VPWR VGND sg13g2_decap_8
XFILLER_40_341 VPWR VGND sg13g2_decap_8
XFILLER_13_599 VPWR VGND sg13g2_decap_8
XFILLER_5_732 VPWR VGND sg13g2_decap_8
XFILLER_4_242 VPWR VGND sg13g2_decap_8
XFILLER_49_931 VPWR VGND sg13g2_decap_8
XFILLER_48_441 VPWR VGND sg13g2_decap_8
XFILLER_24_809 VPWR VGND sg13g2_decap_8
XFILLER_35_124 VPWR VGND sg13g2_decap_8
XFILLER_36_669 VPWR VGND sg13g2_decap_8
XFILLER_17_861 VPWR VGND sg13g2_decap_8
XFILLER_23_319 VPWR VGND sg13g2_decap_8
XFILLER_44_691 VPWR VGND sg13g2_decap_8
XFILLER_32_831 VPWR VGND sg13g2_decap_8
XFILLER_31_330 VPWR VGND sg13g2_decap_8
XFILLER_8_592 VPWR VGND sg13g2_decap_8
XFILLER_6_60 VPWR VGND sg13g2_decap_8
XFILLER_39_452 VPWR VGND sg13g2_decap_8
XFILLER_26_102 VPWR VGND sg13g2_decap_8
XFILLER_27_658 VPWR VGND sg13g2_decap_8
XFILLER_42_628 VPWR VGND sg13g2_decap_8
XFILLER_25_25 VPWR VGND sg13g2_decap_8
XFILLER_26_179 VPWR VGND sg13g2_decap_8
XFILLER_41_116 VPWR VGND sg13g2_decap_8
XFILLER_22_341 VPWR VGND sg13g2_fill_2
XFILLER_23_886 VPWR VGND sg13g2_decap_8
XFILLER_10_536 VPWR VGND sg13g2_decap_8
XFILLER_41_46 VPWR VGND sg13g2_decap_8
XFILLER_6_529 VPWR VGND sg13g2_decap_8
XFILLER_9_4 VPWR VGND sg13g2_decap_8
XFILLER_2_746 VPWR VGND sg13g2_decap_8
XFILLER_1_245 VPWR VGND sg13g2_decap_8
XFILLER_49_238 VPWR VGND sg13g2_decap_8
XFILLER_2_18 VPWR VGND sg13g2_decap_8
XFILLER_46_945 VPWR VGND sg13g2_decap_8
XFILLER_45_411 VPWR VGND sg13g2_decap_8
XFILLER_18_669 VPWR VGND sg13g2_decap_8
XFILLER_45_488 VPWR VGND sg13g2_decap_8
XFILLER_17_168 VPWR VGND sg13g2_decap_8
XFILLER_33_628 VPWR VGND sg13g2_decap_8
XFILLER_32_138 VPWR VGND sg13g2_decap_8
XFILLER_14_864 VPWR VGND sg13g2_decap_8
XFILLER_9_312 VPWR VGND sg13g2_decap_8
XFILLER_13_396 VPWR VGND sg13g2_decap_8
XFILLER_40_193 VPWR VGND sg13g2_decap_8
XFILLER_9_389 VPWR VGND sg13g2_decap_8
XFILLER_37_923 VPWR VGND sg13g2_decap_8
XFILLER_24_606 VPWR VGND sg13g2_decap_8
XFILLER_36_466 VPWR VGND sg13g2_decap_8
XFILLER_23_116 VPWR VGND sg13g2_decap_8
XFILLER_20_845 VPWR VGND sg13g2_decap_8
XFILLER_28_967 VPWR VGND sg13g2_decap_8
XFILLER_43_915 VPWR VGND sg13g2_decap_8
XFILLER_27_455 VPWR VGND sg13g2_decap_8
XFILLER_36_68 VPWR VGND sg13g2_decap_8
XFILLER_42_425 VPWR VGND sg13g2_decap_8
XFILLER_14_116 VPWR VGND sg13g2_decap_8
XFILLER_11_823 VPWR VGND sg13g2_decap_8
XFILLER_23_683 VPWR VGND sg13g2_decap_8
XFILLER_35_1025 VPWR VGND sg13g2_decap_4
XFILLER_10_333 VPWR VGND sg13g2_decap_8
XFILLER_7_805 VPWR VGND sg13g2_decap_8
XFILLER_6_326 VPWR VGND sg13g2_decap_8
XFILLER_2_543 VPWR VGND sg13g2_decap_8
XFILLER_19_923 VPWR VGND sg13g2_decap_8
XFILLER_37_208 VPWR VGND sg13g2_decap_8
XFILLER_46_742 VPWR VGND sg13g2_decap_8
XFILLER_18_466 VPWR VGND sg13g2_decap_8
XFILLER_33_403 VPWR VGND sg13g2_fill_2
XFILLER_45_285 VPWR VGND sg13g2_decap_8
XFILLER_33_425 VPWR VGND sg13g2_decap_8
XFILLER_34_937 VPWR VGND sg13g2_decap_8
XFILLER_42_992 VPWR VGND sg13g2_decap_8
XFILLER_14_661 VPWR VGND sg13g2_decap_8
XFILLER_13_193 VPWR VGND sg13g2_decap_8
XFILLER_9_186 VPWR VGND sg13g2_decap_8
XFILLER_6_893 VPWR VGND sg13g2_decap_8
XFILLER_3_1012 VPWR VGND sg13g2_decap_8
XFILLER_37_720 VPWR VGND sg13g2_decap_8
XFILLER_25_915 VPWR VGND sg13g2_decap_8
XFILLER_36_230 VPWR VGND sg13g2_decap_4
XFILLER_37_797 VPWR VGND sg13g2_decap_8
XFILLER_33_992 VPWR VGND sg13g2_decap_8
XFILLER_40_929 VPWR VGND sg13g2_decap_8
XFILLER_20_642 VPWR VGND sg13g2_decap_8
XFILLER_47_539 VPWR VGND sg13g2_decap_8
XFILLER_47_56 VPWR VGND sg13g2_decap_8
XFILLER_27_252 VPWR VGND sg13g2_decap_8
XFILLER_28_764 VPWR VGND sg13g2_decap_8
XFILLER_43_712 VPWR VGND sg13g2_decap_8
XFILLER_16_937 VPWR VGND sg13g2_decap_8
XFILLER_42_222 VPWR VGND sg13g2_decap_8
XFILLER_15_469 VPWR VGND sg13g2_decap_8
XFILLER_31_918 VPWR VGND sg13g2_decap_8
XFILLER_43_789 VPWR VGND sg13g2_decap_8
XFILLER_24_970 VPWR VGND sg13g2_decap_8
XFILLER_42_299 VPWR VGND sg13g2_decap_8
XFILLER_8_39 VPWR VGND sg13g2_decap_8
XFILLER_11_620 VPWR VGND sg13g2_decap_8
XFILLER_23_480 VPWR VGND sg13g2_decap_8
XFILLER_10_130 VPWR VGND sg13g2_decap_8
XFILLER_7_602 VPWR VGND sg13g2_decap_8
XFILLER_6_123 VPWR VGND sg13g2_decap_8
XFILLER_11_697 VPWR VGND sg13g2_decap_8
XFILLER_7_679 VPWR VGND sg13g2_decap_8
XFILLER_12_81 VPWR VGND sg13g2_decap_8
X_085_ _034_ mod1.bpsk_mod.i_out\[2\] _033_ _051_ VPWR VGND sg13g2_nand3_1
XFILLER_3_830 VPWR VGND sg13g2_decap_8
XFILLER_2_340 VPWR VGND sg13g2_decap_8
XFILLER_19_720 VPWR VGND sg13g2_decap_8
XFILLER_18_263 VPWR VGND sg13g2_decap_8
XFILLER_19_797 VPWR VGND sg13g2_decap_8
XFILLER_34_734 VPWR VGND sg13g2_decap_8
XFILLER_33_222 VPWR VGND sg13g2_decap_8
XFILLER_30_940 VPWR VGND sg13g2_decap_8
XFILLER_6_690 VPWR VGND sg13g2_decap_8
XFILLER_25_1013 VPWR VGND sg13g2_decap_8
XFILLER_44_509 VPWR VGND sg13g2_decap_8
XFILLER_25_712 VPWR VGND sg13g2_decap_8
XFILLER_37_594 VPWR VGND sg13g2_decap_8
XFILLER_13_907 VPWR VGND sg13g2_decap_8
XFILLER_24_222 VPWR VGND sg13g2_decap_8
XFILLER_12_417 VPWR VGND sg13g2_decap_8
XFILLER_25_789 VPWR VGND sg13g2_decap_8
XFILLER_40_726 VPWR VGND sg13g2_decap_8
XFILLER_24_299 VPWR VGND sg13g2_decap_8
XFILLER_33_47 VPWR VGND sg13g2_decap_8
XFILLER_21_962 VPWR VGND sg13g2_decap_8
XFILLER_32_1006 VPWR VGND sg13g2_decap_8
XFILLER_4_627 VPWR VGND sg13g2_decap_8
XFILLER_3_137 VPWR VGND sg13g2_decap_8
XFILLER_0_833 VPWR VGND sg13g2_decap_8
XFILLER_48_826 VPWR VGND sg13g2_decap_8
XFILLER_47_336 VPWR VGND sg13g2_decap_8
XFILLER_16_734 VPWR VGND sg13g2_decap_8
XFILLER_28_561 VPWR VGND sg13g2_decap_8
XFILLER_15_233 VPWR VGND sg13g2_decap_8
XFILLER_43_586 VPWR VGND sg13g2_decap_8
XFILLER_31_715 VPWR VGND sg13g2_decap_8
XFILLER_15_288 VPWR VGND sg13g2_decap_8
XFILLER_30_236 VPWR VGND sg13g2_decap_8
XFILLER_8_900 VPWR VGND sg13g2_decap_8
XFILLER_12_984 VPWR VGND sg13g2_decap_8
XFILLER_8_977 VPWR VGND sg13g2_decap_8
XFILLER_7_476 VPWR VGND sg13g2_decap_8
XFILLER_11_494 VPWR VGND sg13g2_decap_8
X_137_ net14 VGND VPWR _011_ Demo1.qam16_bits\[2\] clknet_2_1__leaf_clk sg13g2_dfrbpq_1
X_068_ net6 net7 _041_ VPWR VGND sg13g2_nor2b_2
XFILLER_31_5 VPWR VGND sg13g2_decap_8
XFILLER_24_4 VPWR VGND sg13g2_decap_8
XFILLER_39_837 VPWR VGND sg13g2_decap_8
XFILLER_38_347 VPWR VGND sg13g2_decap_8
XFILLER_0_1015 VPWR VGND sg13g2_decap_8
XFILLER_0_84 VPWR VGND sg13g2_decap_8
XFILLER_19_594 VPWR VGND sg13g2_decap_8
XFILLER_34_531 VPWR VGND sg13g2_decap_8
XFILLER_22_737 VPWR VGND sg13g2_decap_8
XFILLER_9_60 VPWR VGND sg13g2_decap_8
XFILLER_29_303 VPWR VGND sg13g2_decap_8
XFILLER_28_25 VPWR VGND sg13g2_decap_8
XFILLER_29_347 VPWR VGND sg13g2_fill_1
XFILLER_44_306 VPWR VGND sg13g2_decap_8
XFILLER_37_391 VPWR VGND sg13g2_decap_8
XFILLER_44_68 VPWR VGND sg13g2_decap_8
XFILLER_13_704 VPWR VGND sg13g2_decap_8
XFILLER_25_586 VPWR VGND sg13g2_decap_8
XFILLER_12_214 VPWR VGND sg13g2_decap_8
XFILLER_40_523 VPWR VGND sg13g2_decap_8
XFILLER_8_207 VPWR VGND sg13g2_decap_8
XFILLER_5_914 VPWR VGND sg13g2_decap_8
XFILLER_20_291 VPWR VGND sg13g2_decap_8
XFILLER_5_18 VPWR VGND sg13g2_decap_8
XFILLER_4_424 VPWR VGND sg13g2_decap_8
XFILLER_0_630 VPWR VGND sg13g2_decap_8
XFILLER_48_623 VPWR VGND sg13g2_decap_8
XFILLER_47_133 VPWR VGND sg13g2_decap_8
XFILLER_16_531 VPWR VGND sg13g2_decap_8
XFILLER_35_339 VPWR VGND sg13g2_decap_8
XFILLER_44_873 VPWR VGND sg13g2_decap_8
XFILLER_43_383 VPWR VGND sg13g2_decap_8
XFILLER_31_512 VPWR VGND sg13g2_decap_8
XFILLER_15_1001 VPWR VGND sg13g2_decap_8
XFILLER_12_781 VPWR VGND sg13g2_decap_8
XFILLER_31_589 VPWR VGND sg13g2_decap_8
XFILLER_8_774 VPWR VGND sg13g2_decap_8
XFILLER_11_291 VPWR VGND sg13g2_decap_8
XFILLER_7_273 VPWR VGND sg13g2_decap_8
XFILLER_4_991 VPWR VGND sg13g2_decap_8
XFILLER_39_634 VPWR VGND sg13g2_decap_8
XFILLER_38_144 VPWR VGND sg13g2_decap_8
XFILLER_22_534 VPWR VGND sg13g2_decap_8
XFILLER_10_718 VPWR VGND sg13g2_decap_8
XFILLER_30_26 VPWR VGND sg13g2_decap_8
XFILLER_2_928 VPWR VGND sg13g2_decap_8
XFILLER_1_427 VPWR VGND sg13g2_decap_8
XFILLER_39_46 VPWR VGND sg13g2_decap_8
XFILLER_29_133 VPWR VGND sg13g2_decap_8
XFILLER_44_103 VPWR VGND sg13g2_decap_8
XFILLER_26_840 VPWR VGND sg13g2_decap_8
XFILLER_41_810 VPWR VGND sg13g2_decap_8
XFILLER_13_501 VPWR VGND sg13g2_decap_8
XFILLER_38_1023 VPWR VGND sg13g2_decap_4
XFILLER_40_320 VPWR VGND sg13g2_decap_8
XFILLER_41_887 VPWR VGND sg13g2_decap_8
XFILLER_13_578 VPWR VGND sg13g2_decap_8
XFILLER_40_397 VPWR VGND sg13g2_decap_8
XFILLER_5_711 VPWR VGND sg13g2_decap_8
XFILLER_4_221 VPWR VGND sg13g2_decap_8
XFILLER_5_788 VPWR VGND sg13g2_decap_8
XFILLER_4_298 VPWR VGND sg13g2_decap_8
XFILLER_20_81 VPWR VGND sg13g2_decap_8
XFILLER_49_910 VPWR VGND sg13g2_decap_8
XFILLER_45_1027 VPWR VGND sg13g2_fill_2
XFILLER_48_420 VPWR VGND sg13g2_decap_8
XFILLER_1_994 VPWR VGND sg13g2_decap_8
XFILLER_49_987 VPWR VGND sg13g2_decap_8
XFILLER_35_103 VPWR VGND sg13g2_decap_8
XFILLER_48_497 VPWR VGND sg13g2_decap_8
XFILLER_17_840 VPWR VGND sg13g2_decap_8
XFILLER_36_648 VPWR VGND sg13g2_decap_8
XFILLER_44_670 VPWR VGND sg13g2_decap_8
XFILLER_32_810 VPWR VGND sg13g2_decap_8
XFILLER_43_180 VPWR VGND sg13g2_decap_8
XFILLER_31_386 VPWR VGND sg13g2_decap_8
XFILLER_32_887 VPWR VGND sg13g2_decap_8
XFILLER_8_571 VPWR VGND sg13g2_decap_8
XFILLER_39_431 VPWR VGND sg13g2_decap_8
XFILLER_27_637 VPWR VGND sg13g2_decap_8
XFILLER_42_607 VPWR VGND sg13g2_decap_8
XFILLER_26_158 VPWR VGND sg13g2_decap_8
XFILLER_22_320 VPWR VGND sg13g2_decap_8
XFILLER_23_865 VPWR VGND sg13g2_decap_8
XFILLER_34_180 VPWR VGND sg13g2_decap_8
XFILLER_10_515 VPWR VGND sg13g2_decap_8
XFILLER_6_508 VPWR VGND sg13g2_decap_8
XFILLER_41_25 VPWR VGND sg13g2_decap_8
XFILLER_2_725 VPWR VGND sg13g2_decap_8
XFILLER_1_224 VPWR VGND sg13g2_decap_8
XFILLER_49_217 VPWR VGND sg13g2_decap_8
XFILLER_46_924 VPWR VGND sg13g2_decap_8
XFILLER_18_648 VPWR VGND sg13g2_decap_8
XFILLER_45_467 VPWR VGND sg13g2_decap_8
XFILLER_17_147 VPWR VGND sg13g2_decap_8
XFILLER_33_607 VPWR VGND sg13g2_decap_8
XFILLER_32_117 VPWR VGND sg13g2_decap_8
XFILLER_14_843 VPWR VGND sg13g2_decap_8
XFILLER_41_684 VPWR VGND sg13g2_decap_8
XFILLER_13_375 VPWR VGND sg13g2_decap_8
XFILLER_15_81 VPWR VGND sg13g2_decap_8
XFILLER_9_368 VPWR VGND sg13g2_decap_8
XFILLER_40_172 VPWR VGND sg13g2_decap_8
XFILLER_12_1026 VPWR VGND sg13g2_fill_2
XFILLER_5_585 VPWR VGND sg13g2_decap_8
XFILLER_1_791 VPWR VGND sg13g2_decap_8
XFILLER_49_784 VPWR VGND sg13g2_decap_8
XFILLER_37_902 VPWR VGND sg13g2_decap_8
XFILLER_48_294 VPWR VGND sg13g2_decap_8
XFILLER_36_445 VPWR VGND sg13g2_decap_8
XFILLER_37_979 VPWR VGND sg13g2_decap_8
XFILLER_20_824 VPWR VGND sg13g2_decap_8
XFILLER_32_684 VPWR VGND sg13g2_decap_8
XFILLER_31_194 VPWR VGND sg13g2_decap_8
XFILLER_11_39 VPWR VGND sg13g2_decap_8
XFILLER_27_434 VPWR VGND sg13g2_decap_8
XFILLER_28_946 VPWR VGND sg13g2_decap_8
XFILLER_39_283 VPWR VGND sg13g2_decap_8
XFILLER_42_404 VPWR VGND sg13g2_decap_8
XFILLER_36_47 VPWR VGND sg13g2_decap_8
XFILLER_35_1004 VPWR VGND sg13g2_decap_8
XFILLER_11_802 VPWR VGND sg13g2_decap_8
XFILLER_23_662 VPWR VGND sg13g2_decap_8
XFILLER_10_312 VPWR VGND sg13g2_decap_8
XFILLER_22_194 VPWR VGND sg13g2_decap_8
XFILLER_6_305 VPWR VGND sg13g2_decap_8
XFILLER_11_879 VPWR VGND sg13g2_decap_8
XFILLER_10_389 VPWR VGND sg13g2_decap_8
XFILLER_2_522 VPWR VGND sg13g2_decap_8
XFILLER_2_599 VPWR VGND sg13g2_decap_8
XFILLER_19_902 VPWR VGND sg13g2_decap_8
XFILLER_46_721 VPWR VGND sg13g2_decap_8
XFILLER_18_445 VPWR VGND sg13g2_decap_8
XFILLER_19_979 VPWR VGND sg13g2_decap_8
XFILLER_34_916 VPWR VGND sg13g2_decap_8
XFILLER_46_798 VPWR VGND sg13g2_decap_8
XFILLER_45_264 VPWR VGND sg13g2_decap_8
XFILLER_14_640 VPWR VGND sg13g2_decap_8
XFILLER_42_971 VPWR VGND sg13g2_decap_8
XFILLER_20_109 VPWR VGND sg13g2_decap_8
XFILLER_41_481 VPWR VGND sg13g2_decap_8
XFILLER_13_172 VPWR VGND sg13g2_decap_8
XFILLER_9_165 VPWR VGND sg13g2_decap_8
XFILLER_6_872 VPWR VGND sg13g2_decap_8
XFILLER_5_382 VPWR VGND sg13g2_decap_8
XFILLER_3_95 VPWR VGND sg13g2_decap_8
XFILLER_49_581 VPWR VGND sg13g2_decap_8
XFILLER_37_776 VPWR VGND sg13g2_decap_8
XFILLER_36_275 VPWR VGND sg13g2_decap_8
XFILLER_24_459 VPWR VGND sg13g2_decap_8
XFILLER_40_908 VPWR VGND sg13g2_decap_8
XFILLER_11_109 VPWR VGND sg13g2_decap_8
XFILLER_33_971 VPWR VGND sg13g2_decap_8
XFILLER_20_621 VPWR VGND sg13g2_decap_8
XFILLER_32_481 VPWR VGND sg13g2_decap_8
XFILLER_20_698 VPWR VGND sg13g2_decap_8
XFILLER_4_809 VPWR VGND sg13g2_decap_8
XFILLER_3_319 VPWR VGND sg13g2_decap_8
XFILLER_47_518 VPWR VGND sg13g2_decap_8
XFILLER_47_35 VPWR VGND sg13g2_decap_8
XFILLER_28_743 VPWR VGND sg13g2_decap_8
XFILLER_16_916 VPWR VGND sg13g2_decap_8
XFILLER_27_231 VPWR VGND sg13g2_decap_8
XFILLER_42_201 VPWR VGND sg13g2_decap_8
XFILLER_43_768 VPWR VGND sg13g2_decap_8
XFILLER_15_448 VPWR VGND sg13g2_decap_8
XFILLER_42_278 VPWR VGND sg13g2_decap_8
XFILLER_30_429 VPWR VGND sg13g2_decap_8
XFILLER_8_18 VPWR VGND sg13g2_decap_8
XFILLER_11_676 VPWR VGND sg13g2_decap_8
XFILLER_10_186 VPWR VGND sg13g2_decap_8
XFILLER_7_658 VPWR VGND sg13g2_decap_8
XFILLER_6_102 VPWR VGND sg13g2_decap_8
XFILLER_12_60 VPWR VGND sg13g2_decap_8
X_084_ _050_ mod1.i_out_qpsk\[2\] _045_ VPWR VGND sg13g2_nand2_1
XFILLER_6_179 VPWR VGND sg13g2_decap_8
XFILLER_3_886 VPWR VGND sg13g2_decap_8
XFILLER_2_396 VPWR VGND sg13g2_decap_8
XFILLER_19_776 VPWR VGND sg13g2_decap_8
XFILLER_46_595 VPWR VGND sg13g2_decap_8
XFILLER_34_713 VPWR VGND sg13g2_decap_8
XFILLER_22_919 VPWR VGND sg13g2_decap_8
XFILLER_30_996 VPWR VGND sg13g2_decap_8
XFILLER_29_529 VPWR VGND sg13g2_decap_8
XFILLER_17_49 VPWR VGND sg13g2_decap_8
XFILLER_24_201 VPWR VGND sg13g2_decap_8
XFILLER_37_573 VPWR VGND sg13g2_decap_8
XFILLER_25_768 VPWR VGND sg13g2_decap_8
XFILLER_24_278 VPWR VGND sg13g2_decap_8
XFILLER_40_705 VPWR VGND sg13g2_decap_8
XFILLER_21_941 VPWR VGND sg13g2_decap_8
XFILLER_33_26 VPWR VGND sg13g2_decap_8
XFILLER_4_606 VPWR VGND sg13g2_decap_8
XFILLER_20_495 VPWR VGND sg13g2_decap_8
XFILLER_3_116 VPWR VGND sg13g2_decap_8
XFILLER_0_812 VPWR VGND sg13g2_decap_8
XFILLER_48_805 VPWR VGND sg13g2_decap_8
XFILLER_0_889 VPWR VGND sg13g2_decap_8
XFILLER_47_315 VPWR VGND sg13g2_decap_8
XFILLER_28_540 VPWR VGND sg13g2_decap_8
XFILLER_16_713 VPWR VGND sg13g2_decap_8
XFILLER_15_212 VPWR VGND sg13g2_decap_8
XFILLER_43_565 VPWR VGND sg13g2_decap_8
XFILLER_30_215 VPWR VGND sg13g2_decap_8
XFILLER_12_963 VPWR VGND sg13g2_decap_8
XFILLER_8_956 VPWR VGND sg13g2_decap_8
XFILLER_11_473 VPWR VGND sg13g2_decap_8
XFILLER_23_81 VPWR VGND sg13g2_decap_8
XFILLER_7_455 VPWR VGND sg13g2_decap_8
X_136_ net14 VGND VPWR _005_ Demo1.qam16_bits\[1\] clknet_2_3__leaf_clk sg13g2_dfrbpq_1
X_067_ mod1.qam16_mod.i_level\[3\] _040_ _000_ VPWR VGND net2 sg13g2_nand3b_1
XFILLER_3_683 VPWR VGND sg13g2_decap_8
XFILLER_2_193 VPWR VGND sg13g2_decap_8
XFILLER_39_816 VPWR VGND sg13g2_decap_8
XFILLER_38_326 VPWR VGND sg13g2_decap_8
XFILLER_47_882 VPWR VGND sg13g2_decap_8
XFILLER_19_573 VPWR VGND sg13g2_decap_8
XFILLER_34_510 VPWR VGND sg13g2_decap_8
XFILLER_46_392 VPWR VGND sg13g2_decap_8
XFILLER_0_63 VPWR VGND sg13g2_decap_8
XFILLER_22_716 VPWR VGND sg13g2_decap_8
XFILLER_21_204 VPWR VGND sg13g2_decap_8
XFILLER_34_587 VPWR VGND sg13g2_decap_8
XFILLER_30_793 VPWR VGND sg13g2_decap_8
XFILLER_1_609 VPWR VGND sg13g2_decap_8
XFILLER_0_119 VPWR VGND sg13g2_decap_8
XFILLER_37_370 VPWR VGND sg13g2_decap_8
XFILLER_44_47 VPWR VGND sg13g2_decap_8
XFILLER_25_565 VPWR VGND sg13g2_decap_8
XFILLER_40_502 VPWR VGND sg13g2_decap_8
XFILLER_40_579 VPWR VGND sg13g2_decap_8
XFILLER_20_270 VPWR VGND sg13g2_decap_8
XFILLER_4_403 VPWR VGND sg13g2_decap_8
XFILLER_48_602 VPWR VGND sg13g2_decap_8
XFILLER_47_112 VPWR VGND sg13g2_decap_8
XFILLER_0_686 VPWR VGND sg13g2_decap_8
XFILLER_48_679 VPWR VGND sg13g2_decap_8
XFILLER_47_189 VPWR VGND sg13g2_decap_8
XFILLER_35_318 VPWR VGND sg13g2_decap_8
XFILLER_44_852 VPWR VGND sg13g2_decap_8
XFILLER_16_510 VPWR VGND sg13g2_decap_8
XFILLER_18_81 VPWR VGND sg13g2_decap_8
XFILLER_29_893 VPWR VGND sg13g2_decap_8
XFILLER_43_362 VPWR VGND sg13g2_decap_8
XFILLER_16_587 VPWR VGND sg13g2_decap_8
XFILLER_31_568 VPWR VGND sg13g2_decap_8
XFILLER_12_760 VPWR VGND sg13g2_decap_8
XFILLER_8_753 VPWR VGND sg13g2_decap_8
XFILLER_11_270 VPWR VGND sg13g2_decap_8
XFILLER_7_252 VPWR VGND sg13g2_decap_8
X_119_ _031_ _003_ _030_ _001_ VPWR VGND sg13g2_a21o_1
XFILLER_4_970 VPWR VGND sg13g2_decap_8
XFILLER_3_480 VPWR VGND sg13g2_decap_8
XFILLER_39_613 VPWR VGND sg13g2_decap_8
XFILLER_22_1017 VPWR VGND sg13g2_decap_8
XFILLER_22_1028 VPWR VGND sg13g2_fill_1
XFILLER_27_819 VPWR VGND sg13g2_decap_8
XFILLER_38_123 VPWR VGND sg13g2_decap_8
XFILLER_26_329 VPWR VGND sg13g2_decap_8
XFILLER_19_381 VPWR VGND sg13g2_decap_4
XFILLER_35_885 VPWR VGND sg13g2_decap_8
XFILLER_22_513 VPWR VGND sg13g2_decap_8
XFILLER_34_384 VPWR VGND sg13g2_decap_8
XFILLER_14_39 VPWR VGND sg13g2_decap_8
XFILLER_30_590 VPWR VGND sg13g2_decap_8
XFILLER_2_907 VPWR VGND sg13g2_decap_8
XFILLER_1_406 VPWR VGND sg13g2_decap_8
XFILLER_39_25 VPWR VGND sg13g2_decap_8
XFILLER_29_112 VPWR VGND sg13g2_decap_8
XFILLER_45_649 VPWR VGND sg13g2_decap_8
XFILLER_17_329 VPWR VGND sg13g2_decap_8
XFILLER_29_189 VPWR VGND sg13g2_decap_4
XFILLER_44_159 VPWR VGND sg13g2_decap_8
XFILLER_38_1002 VPWR VGND sg13g2_decap_8
XFILLER_26_896 VPWR VGND sg13g2_decap_8
XFILLER_41_866 VPWR VGND sg13g2_decap_8
XFILLER_13_557 VPWR VGND sg13g2_decap_8
XFILLER_25_395 VPWR VGND sg13g2_decap_8
XFILLER_40_376 VPWR VGND sg13g2_decap_8
XFILLER_4_200 VPWR VGND sg13g2_decap_8
XFILLER_5_767 VPWR VGND sg13g2_decap_8
XFILLER_20_60 VPWR VGND sg13g2_decap_8
XFILLER_45_1006 VPWR VGND sg13g2_decap_8
XFILLER_4_277 VPWR VGND sg13g2_decap_8
XFILLER_1_973 VPWR VGND sg13g2_decap_8
XFILLER_49_966 VPWR VGND sg13g2_decap_8
XFILLER_0_483 VPWR VGND sg13g2_decap_8
XFILLER_48_476 VPWR VGND sg13g2_decap_8
XFILLER_29_91 VPWR VGND sg13g2_decap_8
XFILLER_36_627 VPWR VGND sg13g2_decap_8
XFILLER_29_690 VPWR VGND sg13g2_decap_8
XFILLER_35_159 VPWR VGND sg13g2_decap_8
XFILLER_16_384 VPWR VGND sg13g2_decap_8
XFILLER_17_896 VPWR VGND sg13g2_decap_8
XFILLER_32_866 VPWR VGND sg13g2_decap_8
XFILLER_31_365 VPWR VGND sg13g2_decap_8
XFILLER_8_550 VPWR VGND sg13g2_decap_8
XFILLER_6_95 VPWR VGND sg13g2_decap_8
XFILLER_39_410 VPWR VGND sg13g2_decap_8
XFILLER_27_616 VPWR VGND sg13g2_decap_8
XFILLER_39_487 VPWR VGND sg13g2_decap_8
XFILLER_26_137 VPWR VGND sg13g2_decap_8
XFILLER_35_682 VPWR VGND sg13g2_decap_8
XFILLER_22_343 VPWR VGND sg13g2_fill_1
XFILLER_23_844 VPWR VGND sg13g2_decap_8
XFILLER_22_376 VPWR VGND sg13g2_decap_8
XFILLER_22_387 VPWR VGND sg13g2_fill_1
XFILLER_2_704 VPWR VGND sg13g2_decap_8
XFILLER_1_203 VPWR VGND sg13g2_decap_8
XFILLER_46_903 VPWR VGND sg13g2_decap_8
XFILLER_18_627 VPWR VGND sg13g2_decap_8
XFILLER_45_446 VPWR VGND sg13g2_decap_8
XFILLER_17_126 VPWR VGND sg13g2_decap_8
XFILLER_14_822 VPWR VGND sg13g2_decap_8
XFILLER_26_693 VPWR VGND sg13g2_decap_8
XFILLER_41_663 VPWR VGND sg13g2_decap_8
XFILLER_13_354 VPWR VGND sg13g2_decap_8
XFILLER_14_899 VPWR VGND sg13g2_decap_8
XFILLER_15_60 VPWR VGND sg13g2_decap_8
XFILLER_40_151 VPWR VGND sg13g2_decap_8
XFILLER_9_347 VPWR VGND sg13g2_decap_8
XFILLER_12_1005 VPWR VGND sg13g2_decap_8
XFILLER_5_564 VPWR VGND sg13g2_decap_8
XFILLER_49_7 VPWR VGND sg13g2_decap_8
XFILLER_1_770 VPWR VGND sg13g2_decap_8
XFILLER_0_280 VPWR VGND sg13g2_decap_8
XFILLER_49_763 VPWR VGND sg13g2_decap_8
XFILLER_48_273 VPWR VGND sg13g2_decap_8
XFILLER_36_424 VPWR VGND sg13g2_decap_8
XFILLER_37_958 VPWR VGND sg13g2_decap_8
XFILLER_17_693 VPWR VGND sg13g2_decap_8
XFILLER_20_803 VPWR VGND sg13g2_decap_8
XFILLER_32_663 VPWR VGND sg13g2_decap_8
XFILLER_31_173 VPWR VGND sg13g2_decap_8
XFILLER_11_18 VPWR VGND sg13g2_decap_8
XFILLER_28_1023 VPWR VGND sg13g2_decap_4
XFILLER_28_925 VPWR VGND sg13g2_decap_8
XFILLER_27_413 VPWR VGND sg13g2_decap_8
XFILLER_36_26 VPWR VGND sg13g2_decap_8
XFILLER_36_991 VPWR VGND sg13g2_decap_8
XFILLER_23_641 VPWR VGND sg13g2_decap_8
XFILLER_22_151 VPWR VGND sg13g2_decap_8
XFILLER_11_858 VPWR VGND sg13g2_decap_8
XFILLER_22_173 VPWR VGND sg13g2_decap_8
XFILLER_10_368 VPWR VGND sg13g2_decap_8
XFILLER_2_501 VPWR VGND sg13g2_decap_8
XFILLER_2_578 VPWR VGND sg13g2_decap_8
XFILLER_46_700 VPWR VGND sg13g2_decap_8
XFILLER_18_424 VPWR VGND sg13g2_decap_8
XFILLER_19_958 VPWR VGND sg13g2_decap_8
XFILLER_46_777 VPWR VGND sg13g2_decap_8
XFILLER_45_243 VPWR VGND sg13g2_decap_8
XFILLER_27_980 VPWR VGND sg13g2_decap_8
XFILLER_42_950 VPWR VGND sg13g2_decap_8
XFILLER_26_81 VPWR VGND sg13g2_decap_8
XFILLER_26_490 VPWR VGND sg13g2_decap_8
XFILLER_41_460 VPWR VGND sg13g2_decap_8
XFILLER_13_151 VPWR VGND sg13g2_decap_8
XFILLER_14_696 VPWR VGND sg13g2_decap_8
XFILLER_9_144 VPWR VGND sg13g2_decap_8
XFILLER_6_851 VPWR VGND sg13g2_decap_8
XFILLER_5_361 VPWR VGND sg13g2_decap_8
XFILLER_3_74 VPWR VGND sg13g2_decap_8
XFILLER_49_560 VPWR VGND sg13g2_decap_8
XFILLER_37_755 VPWR VGND sg13g2_decap_8
XFILLER_18_991 VPWR VGND sg13g2_decap_8
XFILLER_36_254 VPWR VGND sg13g2_decap_8
XFILLER_17_490 VPWR VGND sg13g2_decap_8
XFILLER_24_438 VPWR VGND sg13g2_decap_8
XFILLER_33_950 VPWR VGND sg13g2_decap_8
XFILLER_20_600 VPWR VGND sg13g2_decap_8
XFILLER_32_460 VPWR VGND sg13g2_decap_8
XFILLER_22_39 VPWR VGND sg13g2_decap_8
XFILLER_20_677 VPWR VGND sg13g2_decap_8
XFILLER_47_14 VPWR VGND sg13g2_decap_8
XFILLER_41_1020 VPWR VGND sg13g2_decap_8
XFILLER_27_210 VPWR VGND sg13g2_decap_8
XFILLER_28_722 VPWR VGND sg13g2_decap_8
XFILLER_15_427 VPWR VGND sg13g2_decap_8
XFILLER_28_799 VPWR VGND sg13g2_decap_8
XFILLER_43_747 VPWR VGND sg13g2_decap_8
XFILLER_27_287 VPWR VGND sg13g2_fill_1
XFILLER_42_257 VPWR VGND sg13g2_decap_8
XFILLER_30_408 VPWR VGND sg13g2_decap_8
XFILLER_11_655 VPWR VGND sg13g2_decap_8
XFILLER_10_165 VPWR VGND sg13g2_decap_8
XFILLER_7_637 VPWR VGND sg13g2_decap_8
XFILLER_6_158 VPWR VGND sg13g2_decap_8
X_083_ _049_ mod1.i_out_8psk\[2\] _041_ VPWR VGND sg13g2_nand2_1
XFILLER_3_865 VPWR VGND sg13g2_decap_8
XFILLER_2_375 VPWR VGND sg13g2_decap_8
XFILLER_38_519 VPWR VGND sg13g2_decap_8
XFILLER_18_221 VPWR VGND sg13g2_decap_8
XFILLER_19_755 VPWR VGND sg13g2_decap_8
XFILLER_46_574 VPWR VGND sg13g2_decap_8
XFILLER_37_91 VPWR VGND sg13g2_decap_8
XFILLER_18_298 VPWR VGND sg13g2_decap_8
XFILLER_34_769 VPWR VGND sg13g2_decap_8
XFILLER_33_257 VPWR VGND sg13g2_decap_4
XFILLER_33_279 VPWR VGND sg13g2_decap_4
XFILLER_15_994 VPWR VGND sg13g2_decap_8
XFILLER_14_493 VPWR VGND sg13g2_decap_8
XFILLER_30_975 VPWR VGND sg13g2_decap_8
XFILLER_29_508 VPWR VGND sg13g2_decap_8
XFILLER_17_28 VPWR VGND sg13g2_decap_8
XFILLER_37_552 VPWR VGND sg13g2_decap_8
XFILLER_25_747 VPWR VGND sg13g2_decap_8
XFILLER_24_257 VPWR VGND sg13g2_decap_8
XFILLER_21_920 VPWR VGND sg13g2_decap_8
XFILLER_20_474 VPWR VGND sg13g2_decap_8
XFILLER_21_997 VPWR VGND sg13g2_decap_8
XFILLER_0_868 VPWR VGND sg13g2_decap_8
XFILLER_43_544 VPWR VGND sg13g2_decap_8
XFILLER_28_596 VPWR VGND sg13g2_decap_8
XFILLER_16_769 VPWR VGND sg13g2_decap_8
XFILLER_12_942 VPWR VGND sg13g2_decap_8
XFILLER_8_935 VPWR VGND sg13g2_decap_8
XFILLER_11_452 VPWR VGND sg13g2_decap_8
XFILLER_23_60 VPWR VGND sg13g2_decap_8
XFILLER_7_434 VPWR VGND sg13g2_decap_8
X_135_ net14 VGND VPWR _004_ Demo1.qam16_bits\[0\] clknet_2_1__leaf_clk sg13g2_dfrbpq_1
X_066_ net3 net4 _040_ VPWR VGND sg13g2_nor2_2
XFILLER_48_1015 VPWR VGND sg13g2_decap_8
XFILLER_3_662 VPWR VGND sg13g2_decap_8
XFILLER_2_172 VPWR VGND sg13g2_decap_8
XFILLER_38_305 VPWR VGND sg13g2_decap_8
XFILLER_47_861 VPWR VGND sg13g2_decap_8
XFILLER_0_42 VPWR VGND sg13g2_decap_8
XFILLER_19_552 VPWR VGND sg13g2_decap_8
XFILLER_46_371 VPWR VGND sg13g2_decap_8
XFILLER_34_566 VPWR VGND sg13g2_decap_8
XFILLER_15_791 VPWR VGND sg13g2_decap_8
XFILLER_14_290 VPWR VGND sg13g2_decap_8
XFILLER_21_249 VPWR VGND sg13g2_decap_8
XFILLER_9_95 VPWR VGND sg13g2_decap_8
XFILLER_30_772 VPWR VGND sg13g2_decap_8
XFILLER_29_338 VPWR VGND sg13g2_decap_8
XFILLER_38_883 VPWR VGND sg13g2_decap_8
XFILLER_44_26 VPWR VGND sg13g2_decap_8
XFILLER_25_544 VPWR VGND sg13g2_decap_8
XFILLER_13_739 VPWR VGND sg13g2_decap_8
XFILLER_12_249 VPWR VGND sg13g2_decap_8
XFILLER_40_558 VPWR VGND sg13g2_decap_8
XFILLER_21_794 VPWR VGND sg13g2_decap_8
XFILLER_5_949 VPWR VGND sg13g2_decap_8
XFILLER_4_459 VPWR VGND sg13g2_decap_8
XFILLER_0_665 VPWR VGND sg13g2_decap_8
XFILLER_48_658 VPWR VGND sg13g2_decap_8
XFILLER_36_809 VPWR VGND sg13g2_decap_8
XFILLER_47_168 VPWR VGND sg13g2_decap_8
XFILLER_18_60 VPWR VGND sg13g2_decap_8
XFILLER_29_872 VPWR VGND sg13g2_decap_8
XFILLER_44_831 VPWR VGND sg13g2_decap_8
XFILLER_28_382 VPWR VGND sg13g2_decap_8
XFILLER_43_341 VPWR VGND sg13g2_decap_8
XFILLER_16_566 VPWR VGND sg13g2_decap_8
XFILLER_31_547 VPWR VGND sg13g2_decap_8
XFILLER_8_732 VPWR VGND sg13g2_decap_8
XFILLER_7_231 VPWR VGND sg13g2_decap_8
X_118_ net9 net8 _037_ _031_ VPWR VGND sg13g2_nor3_1
XFILLER_38_102 VPWR VGND sg13g2_decap_8
XFILLER_39_669 VPWR VGND sg13g2_decap_8
XFILLER_26_308 VPWR VGND sg13g2_fill_1
XFILLER_38_179 VPWR VGND sg13g2_decap_8
XFILLER_19_360 VPWR VGND sg13g2_decap_8
XFILLER_34_352 VPWR VGND sg13g2_decap_4
XFILLER_35_864 VPWR VGND sg13g2_decap_8
XFILLER_14_18 VPWR VGND sg13g2_decap_8
XFILLER_22_569 VPWR VGND sg13g2_decap_8
XFILLER_18_809 VPWR VGND sg13g2_decap_8
XFILLER_45_628 VPWR VGND sg13g2_decap_8
XFILLER_17_308 VPWR VGND sg13g2_decap_8
XFILLER_29_168 VPWR VGND sg13g2_decap_8
XFILLER_44_138 VPWR VGND sg13g2_decap_8
XFILLER_38_680 VPWR VGND sg13g2_decap_8
XFILLER_26_875 VPWR VGND sg13g2_decap_8
XFILLER_25_374 VPWR VGND sg13g2_decap_8
XFILLER_41_845 VPWR VGND sg13g2_decap_8
XFILLER_13_536 VPWR VGND sg13g2_decap_8
XFILLER_9_529 VPWR VGND sg13g2_decap_8
XFILLER_40_355 VPWR VGND sg13g2_decap_8
XFILLER_21_591 VPWR VGND sg13g2_decap_8
XFILLER_5_746 VPWR VGND sg13g2_decap_8
XFILLER_4_256 VPWR VGND sg13g2_decap_8
XFILLER_1_952 VPWR VGND sg13g2_decap_8
XFILLER_0_462 VPWR VGND sg13g2_decap_8
XFILLER_49_945 VPWR VGND sg13g2_decap_8
XFILLER_29_70 VPWR VGND sg13g2_decap_8
XFILLER_48_455 VPWR VGND sg13g2_decap_8
XFILLER_36_606 VPWR VGND sg13g2_decap_8
XFILLER_35_138 VPWR VGND sg13g2_decap_8
XFILLER_17_875 VPWR VGND sg13g2_decap_8
XFILLER_28_190 VPWR VGND sg13g2_decap_8
XFILLER_16_363 VPWR VGND sg13g2_decap_8
XFILLER_31_344 VPWR VGND sg13g2_decap_8
XFILLER_32_845 VPWR VGND sg13g2_decap_8
XFILLER_6_74 VPWR VGND sg13g2_decap_8
XFILLER_6_1012 VPWR VGND sg13g2_decap_8
XFILLER_39_466 VPWR VGND sg13g2_decap_8
XFILLER_26_116 VPWR VGND sg13g2_decap_8
XFILLER_23_823 VPWR VGND sg13g2_decap_8
XFILLER_25_39 VPWR VGND sg13g2_decap_8
XFILLER_35_661 VPWR VGND sg13g2_decap_8
XFILLER_22_355 VPWR VGND sg13g2_decap_8
XFILLER_1_259 VPWR VGND sg13g2_decap_8
XFILLER_18_606 VPWR VGND sg13g2_decap_8
XFILLER_46_959 VPWR VGND sg13g2_decap_8
XFILLER_45_425 VPWR VGND sg13g2_decap_8
XFILLER_17_105 VPWR VGND sg13g2_decap_8
XFILLER_14_801 VPWR VGND sg13g2_decap_8
XFILLER_26_672 VPWR VGND sg13g2_decap_8
XFILLER_41_642 VPWR VGND sg13g2_decap_8
XFILLER_13_333 VPWR VGND sg13g2_decap_8
XFILLER_25_182 VPWR VGND sg13g2_decap_8
XFILLER_14_878 VPWR VGND sg13g2_decap_8
XFILLER_40_130 VPWR VGND sg13g2_decap_8
XFILLER_9_326 VPWR VGND sg13g2_decap_8
XFILLER_12_1028 VPWR VGND sg13g2_fill_1
XFILLER_5_543 VPWR VGND sg13g2_decap_8
XFILLER_31_82 VPWR VGND sg13g2_decap_8
XFILLER_49_742 VPWR VGND sg13g2_decap_8
XFILLER_48_252 VPWR VGND sg13g2_decap_8
XFILLER_36_403 VPWR VGND sg13g2_decap_8
XFILLER_37_937 VPWR VGND sg13g2_decap_8
XFILLER_45_992 VPWR VGND sg13g2_decap_8
XFILLER_17_672 VPWR VGND sg13g2_decap_8
XFILLER_16_193 VPWR VGND sg13g2_decap_8
XFILLER_32_642 VPWR VGND sg13g2_decap_8
XFILLER_31_152 VPWR VGND sg13g2_decap_8
XFILLER_20_859 VPWR VGND sg13g2_decap_8
XFILLER_9_893 VPWR VGND sg13g2_decap_8
XFILLER_28_1002 VPWR VGND sg13g2_decap_8
XFILLER_28_904 VPWR VGND sg13g2_decap_8
XFILLER_39_263 VPWR VGND sg13g2_decap_8
XFILLER_15_609 VPWR VGND sg13g2_decap_8
XFILLER_27_469 VPWR VGND sg13g2_decap_8
XFILLER_43_929 VPWR VGND sg13g2_decap_8
XFILLER_36_970 VPWR VGND sg13g2_decap_8
XFILLER_42_439 VPWR VGND sg13g2_decap_8
XFILLER_23_620 VPWR VGND sg13g2_decap_8
XFILLER_22_130 VPWR VGND sg13g2_decap_8
XFILLER_11_837 VPWR VGND sg13g2_decap_8
XFILLER_23_697 VPWR VGND sg13g2_decap_8
XFILLER_10_347 VPWR VGND sg13g2_decap_8
XFILLER_7_819 VPWR VGND sg13g2_decap_8
XFILLER_2_557 VPWR VGND sg13g2_decap_8
XFILLER_18_403 VPWR VGND sg13g2_decap_8
XFILLER_19_937 VPWR VGND sg13g2_decap_8
XFILLER_46_756 VPWR VGND sg13g2_decap_8
XFILLER_45_222 VPWR VGND sg13g2_decap_8
XFILLER_26_60 VPWR VGND sg13g2_decap_8
XFILLER_45_299 VPWR VGND sg13g2_decap_8
XFILLER_33_439 VPWR VGND sg13g2_decap_8
XFILLER_13_130 VPWR VGND sg13g2_decap_8
XFILLER_14_675 VPWR VGND sg13g2_decap_8
XFILLER_9_123 VPWR VGND sg13g2_decap_8
XFILLER_6_830 VPWR VGND sg13g2_decap_8
XFILLER_5_340 VPWR VGND sg13g2_decap_8
XFILLER_3_53 VPWR VGND sg13g2_decap_8
XFILLER_3_1026 VPWR VGND sg13g2_fill_2
XFILLER_37_734 VPWR VGND sg13g2_decap_8
XFILLER_36_222 VPWR VGND sg13g2_fill_1
XFILLER_18_970 VPWR VGND sg13g2_decap_8
XFILLER_25_929 VPWR VGND sg13g2_decap_8
XFILLER_20_656 VPWR VGND sg13g2_decap_8
XFILLER_22_18 VPWR VGND sg13g2_decap_8
XFILLER_9_690 VPWR VGND sg13g2_decap_8
XFILLER_28_701 VPWR VGND sg13g2_decap_8
XFILLER_43_726 VPWR VGND sg13g2_decap_8
XFILLER_15_406 VPWR VGND sg13g2_decap_8
XFILLER_27_266 VPWR VGND sg13g2_decap_8
XFILLER_28_778 VPWR VGND sg13g2_decap_8
XFILLER_42_236 VPWR VGND sg13g2_decap_8
XFILLER_24_984 VPWR VGND sg13g2_decap_8
XFILLER_7_616 VPWR VGND sg13g2_decap_8
XFILLER_11_634 VPWR VGND sg13g2_decap_8
XFILLER_23_494 VPWR VGND sg13g2_decap_8
XFILLER_10_144 VPWR VGND sg13g2_decap_8
XFILLER_6_137 VPWR VGND sg13g2_decap_8
X_082_ VGND VPWR _048_ net26 _047_ _046_ sg13g2_a21oi_2
XFILLER_12_95 VPWR VGND sg13g2_decap_8
XFILLER_3_844 VPWR VGND sg13g2_decap_8
XFILLER_2_354 VPWR VGND sg13g2_decap_8
XFILLER_18_200 VPWR VGND sg13g2_decap_8
XFILLER_19_734 VPWR VGND sg13g2_decap_8
XFILLER_46_553 VPWR VGND sg13g2_decap_8
XFILLER_18_277 VPWR VGND sg13g2_decap_8
XFILLER_33_203 VPWR VGND sg13g2_decap_8
XFILLER_37_70 VPWR VGND sg13g2_decap_8
XFILLER_33_236 VPWR VGND sg13g2_decap_8
XFILLER_34_748 VPWR VGND sg13g2_decap_8
XFILLER_15_973 VPWR VGND sg13g2_decap_8
XFILLER_18_1012 VPWR VGND sg13g2_decap_8
XFILLER_21_409 VPWR VGND sg13g2_decap_8
XFILLER_14_472 VPWR VGND sg13g2_decap_8
XFILLER_30_954 VPWR VGND sg13g2_decap_8
XFILLER_25_1027 VPWR VGND sg13g2_fill_2
XFILLER_37_531 VPWR VGND sg13g2_decap_8
XFILLER_25_726 VPWR VGND sg13g2_decap_8
XFILLER_24_236 VPWR VGND sg13g2_decap_8
XFILLER_20_453 VPWR VGND sg13g2_decap_8
XFILLER_21_976 VPWR VGND sg13g2_decap_8
XFILLER_0_847 VPWR VGND sg13g2_decap_8
XFILLER_28_575 VPWR VGND sg13g2_decap_8
XFILLER_43_523 VPWR VGND sg13g2_decap_8
XFILLER_16_748 VPWR VGND sg13g2_decap_8
XFILLER_15_247 VPWR VGND sg13g2_decap_8
XFILLER_12_921 VPWR VGND sg13g2_decap_8
XFILLER_24_781 VPWR VGND sg13g2_decap_8
XFILLER_31_729 VPWR VGND sg13g2_decap_8
XFILLER_8_914 VPWR VGND sg13g2_decap_8
XFILLER_11_431 VPWR VGND sg13g2_decap_8
XFILLER_7_413 VPWR VGND sg13g2_decap_8
XFILLER_12_998 VPWR VGND sg13g2_decap_8
X_134_ net15 VGND VPWR _013_ mod1.i_out_qpsk\[2\] clknet_2_2__leaf_clk sg13g2_dfrbpq_1
X_065_ _039_ _032_ mod1.qam16_mod.i_level\[3\] VPWR VGND sg13g2_nand2_2
XFILLER_3_641 VPWR VGND sg13g2_decap_8
XFILLER_2_151 VPWR VGND sg13g2_decap_8
XFILLER_47_840 VPWR VGND sg13g2_decap_8
XFILLER_48_91 VPWR VGND sg13g2_decap_8
XFILLER_19_531 VPWR VGND sg13g2_decap_8
XFILLER_46_350 VPWR VGND sg13g2_decap_8
XFILLER_0_21 VPWR VGND sg13g2_decap_8
XFILLER_0_98 VPWR VGND sg13g2_decap_8
XFILLER_34_545 VPWR VGND sg13g2_decap_8
XFILLER_15_770 VPWR VGND sg13g2_decap_8
XFILLER_21_228 VPWR VGND sg13g2_decap_8
XFILLER_9_74 VPWR VGND sg13g2_decap_8
XFILLER_30_751 VPWR VGND sg13g2_decap_8
XFILLER_7_980 VPWR VGND sg13g2_decap_8
XFILLER_28_39 VPWR VGND sg13g2_decap_8
XFILLER_29_317 VPWR VGND sg13g2_decap_8
XFILLER_38_862 VPWR VGND sg13g2_decap_8
XFILLER_25_523 VPWR VGND sg13g2_decap_8
XFILLER_13_718 VPWR VGND sg13g2_decap_8
XFILLER_12_228 VPWR VGND sg13g2_decap_8
XFILLER_40_537 VPWR VGND sg13g2_decap_8
XFILLER_21_773 VPWR VGND sg13g2_decap_8
XFILLER_5_928 VPWR VGND sg13g2_decap_8
XFILLER_4_438 VPWR VGND sg13g2_decap_8
XFILLER_0_644 VPWR VGND sg13g2_decap_8
XFILLER_48_637 VPWR VGND sg13g2_decap_8
XFILLER_47_147 VPWR VGND sg13g2_decap_8
XFILLER_29_851 VPWR VGND sg13g2_decap_8
XFILLER_44_810 VPWR VGND sg13g2_decap_8
XFILLER_43_320 VPWR VGND sg13g2_decap_8
XFILLER_16_545 VPWR VGND sg13g2_decap_8
XFILLER_44_887 VPWR VGND sg13g2_decap_8
XFILLER_31_526 VPWR VGND sg13g2_decap_8
XFILLER_43_397 VPWR VGND sg13g2_decap_8
XFILLER_34_82 VPWR VGND sg13g2_decap_8
XFILLER_8_711 VPWR VGND sg13g2_decap_8
XFILLER_15_1015 VPWR VGND sg13g2_decap_8
XFILLER_7_210 VPWR VGND sg13g2_decap_8
XFILLER_12_795 VPWR VGND sg13g2_decap_8
XFILLER_8_788 VPWR VGND sg13g2_decap_8
X_117_ net20 _041_ _003_ VPWR VGND sg13g2_and2_1
XFILLER_7_287 VPWR VGND sg13g2_decap_8
XFILLER_22_4 VPWR VGND sg13g2_decap_8
XFILLER_39_648 VPWR VGND sg13g2_decap_8
XFILLER_38_158 VPWR VGND sg13g2_decap_8
XFILLER_34_331 VPWR VGND sg13g2_decap_8
XFILLER_35_843 VPWR VGND sg13g2_decap_8
XFILLER_22_548 VPWR VGND sg13g2_decap_8
XFILLER_45_607 VPWR VGND sg13g2_decap_8
XFILLER_29_147 VPWR VGND sg13g2_decap_8
XFILLER_44_117 VPWR VGND sg13g2_decap_8
XFILLER_26_854 VPWR VGND sg13g2_decap_8
XFILLER_37_180 VPWR VGND sg13g2_decap_8
XFILLER_41_824 VPWR VGND sg13g2_decap_8
XFILLER_13_515 VPWR VGND sg13g2_decap_8
XFILLER_25_353 VPWR VGND sg13g2_fill_2
XFILLER_9_508 VPWR VGND sg13g2_decap_8
XFILLER_40_334 VPWR VGND sg13g2_decap_8
XFILLER_21_570 VPWR VGND sg13g2_decap_8
XFILLER_5_725 VPWR VGND sg13g2_decap_8
XFILLER_4_235 VPWR VGND sg13g2_decap_8
XFILLER_20_95 VPWR VGND sg13g2_decap_8
XFILLER_1_931 VPWR VGND sg13g2_decap_8
XFILLER_49_924 VPWR VGND sg13g2_decap_8
XFILLER_0_441 VPWR VGND sg13g2_decap_8
XFILLER_48_434 VPWR VGND sg13g2_decap_8
XFILLER_35_117 VPWR VGND sg13g2_decap_8
XFILLER_16_342 VPWR VGND sg13g2_decap_8
XFILLER_17_854 VPWR VGND sg13g2_decap_8
XFILLER_44_684 VPWR VGND sg13g2_decap_8
XFILLER_32_824 VPWR VGND sg13g2_decap_8
XFILLER_43_194 VPWR VGND sg13g2_decap_8
XFILLER_31_323 VPWR VGND sg13g2_decap_8
XFILLER_12_592 VPWR VGND sg13g2_decap_8
XFILLER_8_585 VPWR VGND sg13g2_decap_8
XFILLER_6_53 VPWR VGND sg13g2_decap_8
XFILLER_39_445 VPWR VGND sg13g2_decap_8
XFILLER_25_18 VPWR VGND sg13g2_decap_8
XFILLER_35_640 VPWR VGND sg13g2_decap_8
XFILLER_23_802 VPWR VGND sg13g2_decap_8
XFILLER_41_109 VPWR VGND sg13g2_decap_8
XFILLER_22_334 VPWR VGND sg13g2_decap_8
XFILLER_34_194 VPWR VGND sg13g2_decap_4
XFILLER_23_879 VPWR VGND sg13g2_decap_8
XFILLER_10_529 VPWR VGND sg13g2_decap_8
XFILLER_31_890 VPWR VGND sg13g2_decap_8
XFILLER_41_39 VPWR VGND sg13g2_decap_8
XFILLER_2_739 VPWR VGND sg13g2_decap_8
XFILLER_1_238 VPWR VGND sg13g2_decap_8
XFILLER_46_938 VPWR VGND sg13g2_decap_8
XFILLER_45_404 VPWR VGND sg13g2_decap_8
Xheichips25_template_40 VPWR VGND uio_oe[7] sg13g2_tiehi
XFILLER_26_651 VPWR VGND sg13g2_decap_8
XFILLER_41_621 VPWR VGND sg13g2_decap_8
XFILLER_13_312 VPWR VGND sg13g2_decap_8
XFILLER_14_857 VPWR VGND sg13g2_decap_8
XFILLER_25_161 VPWR VGND sg13g2_decap_8
XFILLER_9_305 VPWR VGND sg13g2_decap_8
XFILLER_41_698 VPWR VGND sg13g2_decap_8
XFILLER_13_389 VPWR VGND sg13g2_decap_8
XFILLER_15_95 VPWR VGND sg13g2_decap_8
XFILLER_40_186 VPWR VGND sg13g2_decap_8
XFILLER_5_522 VPWR VGND sg13g2_decap_8
XFILLER_31_61 VPWR VGND sg13g2_decap_8
XFILLER_5_599 VPWR VGND sg13g2_decap_8
XFILLER_49_721 VPWR VGND sg13g2_decap_8
XFILLER_48_231 VPWR VGND sg13g2_decap_8
XFILLER_37_916 VPWR VGND sg13g2_decap_8
XFILLER_49_798 VPWR VGND sg13g2_decap_8
XFILLER_36_459 VPWR VGND sg13g2_decap_8
XFILLER_45_971 VPWR VGND sg13g2_decap_8
XFILLER_17_651 VPWR VGND sg13g2_decap_8
XFILLER_23_109 VPWR VGND sg13g2_decap_8
XFILLER_44_481 VPWR VGND sg13g2_decap_8
XFILLER_16_172 VPWR VGND sg13g2_decap_8
XFILLER_32_621 VPWR VGND sg13g2_decap_8
XFILLER_31_131 VPWR VGND sg13g2_decap_8
XFILLER_20_838 VPWR VGND sg13g2_decap_8
XFILLER_32_698 VPWR VGND sg13g2_decap_8
XFILLER_9_872 VPWR VGND sg13g2_decap_8
XFILLER_8_382 VPWR VGND sg13g2_decap_8
XFILLER_39_242 VPWR VGND sg13g2_decap_8
XFILLER_43_908 VPWR VGND sg13g2_decap_8
XFILLER_27_448 VPWR VGND sg13g2_decap_8
XFILLER_39_297 VPWR VGND sg13g2_decap_8
XFILLER_42_418 VPWR VGND sg13g2_decap_8
XFILLER_14_109 VPWR VGND sg13g2_decap_8
XFILLER_11_816 VPWR VGND sg13g2_decap_8
XFILLER_23_676 VPWR VGND sg13g2_decap_8
XFILLER_35_1018 VPWR VGND sg13g2_decap_8
XFILLER_10_326 VPWR VGND sg13g2_decap_8
XFILLER_6_319 VPWR VGND sg13g2_decap_8
XFILLER_2_536 VPWR VGND sg13g2_decap_8
XFILLER_19_916 VPWR VGND sg13g2_decap_8
XFILLER_46_735 VPWR VGND sg13g2_decap_8
XFILLER_45_201 VPWR VGND sg13g2_decap_8
XFILLER_18_459 VPWR VGND sg13g2_decap_8
XFILLER_45_278 VPWR VGND sg13g2_decap_8
XFILLER_33_418 VPWR VGND sg13g2_decap_8
XFILLER_14_654 VPWR VGND sg13g2_decap_8
XFILLER_42_985 VPWR VGND sg13g2_decap_8
XFILLER_9_102 VPWR VGND sg13g2_decap_8
XFILLER_41_495 VPWR VGND sg13g2_decap_8
XFILLER_13_186 VPWR VGND sg13g2_decap_8
XFILLER_42_82 VPWR VGND sg13g2_decap_8
XFILLER_9_179 VPWR VGND sg13g2_decap_8
XFILLER_10_893 VPWR VGND sg13g2_decap_8
XFILLER_6_886 VPWR VGND sg13g2_decap_8
XFILLER_5_396 VPWR VGND sg13g2_decap_8
XFILLER_3_32 VPWR VGND sg13g2_decap_8
XFILLER_3_1005 VPWR VGND sg13g2_decap_8
XFILLER_36_201 VPWR VGND sg13g2_decap_8
XFILLER_37_713 VPWR VGND sg13g2_decap_8
XFILLER_49_595 VPWR VGND sg13g2_decap_8
XFILLER_25_908 VPWR VGND sg13g2_decap_8
XFILLER_36_234 VPWR VGND sg13g2_fill_1
XFILLER_33_985 VPWR VGND sg13g2_decap_8
XFILLER_20_635 VPWR VGND sg13g2_decap_8
XFILLER_32_495 VPWR VGND sg13g2_decap_8
XFILLER_47_49 VPWR VGND sg13g2_decap_8
XFILLER_28_757 VPWR VGND sg13g2_decap_8
XFILLER_43_705 VPWR VGND sg13g2_decap_8
XFILLER_27_245 VPWR VGND sg13g2_decap_8
XFILLER_42_215 VPWR VGND sg13g2_decap_8
XFILLER_24_963 VPWR VGND sg13g2_decap_8
XFILLER_11_613 VPWR VGND sg13g2_decap_8
XFILLER_23_473 VPWR VGND sg13g2_decap_8
XFILLER_10_123 VPWR VGND sg13g2_decap_8
XFILLER_6_116 VPWR VGND sg13g2_decap_8
X_081_ net7 net6 Demo1.qam16_bits\[3\] _048_ VPWR VGND sg13g2_nor3_1
XFILLER_12_74 VPWR VGND sg13g2_decap_8
XFILLER_3_823 VPWR VGND sg13g2_decap_8
XFILLER_2_333 VPWR VGND sg13g2_decap_8
XFILLER_19_713 VPWR VGND sg13g2_decap_8
XFILLER_46_532 VPWR VGND sg13g2_decap_8
XFILLER_18_256 VPWR VGND sg13g2_decap_8
XFILLER_34_727 VPWR VGND sg13g2_decap_8
XFILLER_15_952 VPWR VGND sg13g2_decap_8
XFILLER_42_782 VPWR VGND sg13g2_decap_8
XFILLER_14_451 VPWR VGND sg13g2_decap_8
XFILLER_30_933 VPWR VGND sg13g2_decap_8
XFILLER_41_292 VPWR VGND sg13g2_decap_8
XFILLER_41_270 VPWR VGND sg13g2_decap_8
XFILLER_10_690 VPWR VGND sg13g2_decap_8
XFILLER_6_683 VPWR VGND sg13g2_decap_8
XFILLER_5_193 VPWR VGND sg13g2_decap_8
XFILLER_25_1006 VPWR VGND sg13g2_decap_8
XFILLER_49_392 VPWR VGND sg13g2_decap_8
XFILLER_37_510 VPWR VGND sg13g2_decap_8
XFILLER_25_705 VPWR VGND sg13g2_decap_8
XFILLER_24_215 VPWR VGND sg13g2_decap_8
XFILLER_37_587 VPWR VGND sg13g2_decap_8
XFILLER_40_719 VPWR VGND sg13g2_decap_8
XFILLER_33_782 VPWR VGND sg13g2_decap_8
XFILLER_20_432 VPWR VGND sg13g2_decap_8
XFILLER_21_955 VPWR VGND sg13g2_decap_8
XFILLER_32_292 VPWR VGND sg13g2_decap_8
XFILLER_0_826 VPWR VGND sg13g2_decap_8
XFILLER_48_819 VPWR VGND sg13g2_decap_8
XFILLER_47_329 VPWR VGND sg13g2_decap_8
XFILLER_43_502 VPWR VGND sg13g2_decap_8
XFILLER_28_554 VPWR VGND sg13g2_decap_8
XFILLER_15_226 VPWR VGND sg13g2_decap_8
XFILLER_16_727 VPWR VGND sg13g2_decap_8
XFILLER_31_708 VPWR VGND sg13g2_decap_8
XFILLER_43_579 VPWR VGND sg13g2_decap_8
XFILLER_12_900 VPWR VGND sg13g2_decap_8
XFILLER_24_760 VPWR VGND sg13g2_decap_8
XFILLER_11_410 VPWR VGND sg13g2_decap_8
XFILLER_23_281 VPWR VGND sg13g2_decap_8
XFILLER_30_229 VPWR VGND sg13g2_decap_8
XFILLER_12_977 VPWR VGND sg13g2_decap_8
XFILLER_11_487 VPWR VGND sg13g2_decap_8
X_133_ net13 VGND VPWR _012_ mod1.i_out_qpsk\[1\] clknet_2_2__leaf_clk sg13g2_dfrbpq_1
XFILLER_23_95 VPWR VGND sg13g2_decap_8
XFILLER_7_469 VPWR VGND sg13g2_decap_8
X_064_ net12 VPWR _011_ VGND _037_ _038_ sg13g2_o21ai_1
XFILLER_3_620 VPWR VGND sg13g2_decap_8
XFILLER_2_130 VPWR VGND sg13g2_decap_8
XFILLER_3_697 VPWR VGND sg13g2_decap_8
XFILLER_48_70 VPWR VGND sg13g2_decap_8
XFILLER_17_7 VPWR VGND sg13g2_decap_8
XFILLER_19_510 VPWR VGND sg13g2_decap_8
XFILLER_0_1008 VPWR VGND sg13g2_decap_8
XFILLER_47_896 VPWR VGND sg13g2_decap_8
XFILLER_0_77 VPWR VGND sg13g2_decap_8
XFILLER_19_587 VPWR VGND sg13g2_decap_8
XFILLER_34_524 VPWR VGND sg13g2_decap_8
XFILLER_21_218 VPWR VGND sg13g2_decap_4
XFILLER_9_53 VPWR VGND sg13g2_decap_8
XFILLER_30_730 VPWR VGND sg13g2_decap_8
XFILLER_6_480 VPWR VGND sg13g2_decap_8
XFILLER_28_18 VPWR VGND sg13g2_decap_8
XFILLER_38_841 VPWR VGND sg13g2_decap_8
XFILLER_25_502 VPWR VGND sg13g2_decap_8
XFILLER_37_384 VPWR VGND sg13g2_decap_8
XFILLER_12_207 VPWR VGND sg13g2_decap_8
XFILLER_25_579 VPWR VGND sg13g2_decap_8
XFILLER_40_516 VPWR VGND sg13g2_decap_8
XFILLER_21_752 VPWR VGND sg13g2_decap_8
XFILLER_20_284 VPWR VGND sg13g2_decap_8
XFILLER_5_907 VPWR VGND sg13g2_decap_8
XFILLER_4_417 VPWR VGND sg13g2_decap_8
XFILLER_0_623 VPWR VGND sg13g2_decap_8
XFILLER_48_616 VPWR VGND sg13g2_decap_8
XFILLER_47_126 VPWR VGND sg13g2_decap_8
XFILLER_29_830 VPWR VGND sg13g2_decap_8
XFILLER_16_524 VPWR VGND sg13g2_decap_8
XFILLER_18_95 VPWR VGND sg13g2_decap_8
XFILLER_44_866 VPWR VGND sg13g2_decap_8
XFILLER_43_376 VPWR VGND sg13g2_decap_8
XFILLER_31_505 VPWR VGND sg13g2_decap_8
XFILLER_34_61 VPWR VGND sg13g2_decap_8
XFILLER_12_774 VPWR VGND sg13g2_decap_8
XFILLER_11_284 VPWR VGND sg13g2_decap_8
XFILLER_8_767 VPWR VGND sg13g2_decap_8
XFILLER_7_266 VPWR VGND sg13g2_decap_8
X_116_ _033_ net6 net20 _029_ _030_ VPWR VGND sg13g2_nor4_1
XFILLER_4_984 VPWR VGND sg13g2_decap_8
XFILLER_3_494 VPWR VGND sg13g2_decap_8
XFILLER_39_627 VPWR VGND sg13g2_decap_8
XFILLER_15_4 VPWR VGND sg13g2_decap_8
XFILLER_38_137 VPWR VGND sg13g2_decap_8
XFILLER_47_693 VPWR VGND sg13g2_decap_8
XFILLER_34_310 VPWR VGND sg13g2_decap_8
XFILLER_35_822 VPWR VGND sg13g2_decap_8
XFILLER_35_899 VPWR VGND sg13g2_decap_8
XFILLER_22_527 VPWR VGND sg13g2_decap_8
XFILLER_34_398 VPWR VGND sg13g2_decap_8
XFILLER_30_19 VPWR VGND sg13g2_decap_8
XFILLER_39_39 VPWR VGND sg13g2_decap_8
XFILLER_29_126 VPWR VGND sg13g2_decap_8
XFILLER_26_833 VPWR VGND sg13g2_decap_8
XFILLER_25_332 VPWR VGND sg13g2_decap_8
XFILLER_41_803 VPWR VGND sg13g2_decap_8
XFILLER_38_1016 VPWR VGND sg13g2_decap_8
XFILLER_38_1027 VPWR VGND sg13g2_fill_2
XFILLER_40_313 VPWR VGND sg13g2_decap_8
XFILLER_5_704 VPWR VGND sg13g2_decap_8
XFILLER_4_214 VPWR VGND sg13g2_decap_8
XFILLER_1_910 VPWR VGND sg13g2_decap_8
XFILLER_20_74 VPWR VGND sg13g2_decap_8
XFILLER_0_420 VPWR VGND sg13g2_decap_8
XFILLER_49_903 VPWR VGND sg13g2_decap_8
XFILLER_1_987 VPWR VGND sg13g2_decap_8
XFILLER_48_413 VPWR VGND sg13g2_decap_8
XFILLER_0_497 VPWR VGND sg13g2_decap_8
XFILLER_17_833 VPWR VGND sg13g2_decap_8
XFILLER_45_82 VPWR VGND sg13g2_decap_8
XFILLER_44_663 VPWR VGND sg13g2_decap_8
XFILLER_32_803 VPWR VGND sg13g2_decap_8
XFILLER_43_173 VPWR VGND sg13g2_decap_8
XFILLER_16_398 VPWR VGND sg13g2_decap_8
XFILLER_12_571 VPWR VGND sg13g2_decap_8
XFILLER_31_379 VPWR VGND sg13g2_decap_8
XFILLER_40_880 VPWR VGND sg13g2_decap_8
XFILLER_8_564 VPWR VGND sg13g2_decap_8
XFILLER_6_32 VPWR VGND sg13g2_decap_8
XFILLER_4_781 VPWR VGND sg13g2_decap_8
XFILLER_3_291 VPWR VGND sg13g2_decap_8
XFILLER_39_424 VPWR VGND sg13g2_decap_8
XFILLER_48_980 VPWR VGND sg13g2_decap_8
XFILLER_47_490 VPWR VGND sg13g2_decap_8
XFILLER_19_181 VPWR VGND sg13g2_fill_2
XFILLER_19_192 VPWR VGND sg13g2_decap_8
XFILLER_22_313 VPWR VGND sg13g2_decap_8
XFILLER_23_858 VPWR VGND sg13g2_decap_8
XFILLER_34_173 VPWR VGND sg13g2_decap_8
XFILLER_35_696 VPWR VGND sg13g2_decap_8
XFILLER_10_508 VPWR VGND sg13g2_decap_8
XFILLER_41_18 VPWR VGND sg13g2_decap_8
XFILLER_2_718 VPWR VGND sg13g2_decap_8
XFILLER_1_217 VPWR VGND sg13g2_decap_8
XFILLER_44_1020 VPWR VGND sg13g2_decap_8
XFILLER_46_917 VPWR VGND sg13g2_decap_8
Xheichips25_template_30 VPWR VGND uio_out[6] sg13g2_tielo
XFILLER_39_991 VPWR VGND sg13g2_decap_8
XFILLER_26_630 VPWR VGND sg13g2_decap_8
XFILLER_41_600 VPWR VGND sg13g2_decap_8
XFILLER_25_151 VPWR VGND sg13g2_fill_2
XFILLER_14_836 VPWR VGND sg13g2_decap_8
XFILLER_41_677 VPWR VGND sg13g2_decap_8
XFILLER_13_368 VPWR VGND sg13g2_decap_8
XFILLER_15_74 VPWR VGND sg13g2_decap_8
XFILLER_40_165 VPWR VGND sg13g2_decap_8
XFILLER_22_891 VPWR VGND sg13g2_decap_8
XFILLER_5_501 VPWR VGND sg13g2_decap_8
XFILLER_12_1019 VPWR VGND sg13g2_decap_8
XFILLER_31_40 VPWR VGND sg13g2_decap_8
XFILLER_5_578 VPWR VGND sg13g2_decap_8
XFILLER_49_700 VPWR VGND sg13g2_decap_8
XFILLER_48_210 VPWR VGND sg13g2_decap_8
XFILLER_1_784 VPWR VGND sg13g2_decap_8
XFILLER_49_777 VPWR VGND sg13g2_decap_8
XFILLER_0_294 VPWR VGND sg13g2_decap_8
XFILLER_48_287 VPWR VGND sg13g2_decap_8
XFILLER_45_950 VPWR VGND sg13g2_decap_8
XFILLER_17_630 VPWR VGND sg13g2_decap_8
XFILLER_36_438 VPWR VGND sg13g2_decap_8
XFILLER_32_600 VPWR VGND sg13g2_decap_8
XFILLER_44_460 VPWR VGND sg13g2_decap_8
XFILLER_16_151 VPWR VGND sg13g2_decap_8
XFILLER_31_110 VPWR VGND sg13g2_decap_8
XFILLER_20_817 VPWR VGND sg13g2_decap_8
XFILLER_32_677 VPWR VGND sg13g2_decap_8
XFILLER_9_851 VPWR VGND sg13g2_decap_8
XFILLER_31_187 VPWR VGND sg13g2_decap_8
XFILLER_8_361 VPWR VGND sg13g2_decap_8
XFILLER_39_221 VPWR VGND sg13g2_decap_8
XFILLER_28_939 VPWR VGND sg13g2_decap_8
XFILLER_27_427 VPWR VGND sg13g2_decap_8
XFILLER_35_493 VPWR VGND sg13g2_decap_8
XFILLER_23_655 VPWR VGND sg13g2_decap_8
XFILLER_10_305 VPWR VGND sg13g2_decap_8
XFILLER_22_187 VPWR VGND sg13g2_decap_8
XFILLER_2_515 VPWR VGND sg13g2_decap_8
XFILLER_46_714 VPWR VGND sg13g2_decap_8
XFILLER_18_438 VPWR VGND sg13g2_decap_8
XFILLER_34_909 VPWR VGND sg13g2_decap_8
XFILLER_45_257 VPWR VGND sg13g2_decap_8
XFILLER_27_994 VPWR VGND sg13g2_decap_8
XFILLER_42_964 VPWR VGND sg13g2_decap_8
XFILLER_14_633 VPWR VGND sg13g2_decap_8
XFILLER_26_95 VPWR VGND sg13g2_decap_8
XFILLER_41_474 VPWR VGND sg13g2_decap_8
XFILLER_13_165 VPWR VGND sg13g2_decap_8
XFILLER_42_61 VPWR VGND sg13g2_decap_8
XFILLER_9_158 VPWR VGND sg13g2_decap_8
XFILLER_10_872 VPWR VGND sg13g2_decap_8
XFILLER_6_865 VPWR VGND sg13g2_decap_8
XFILLER_47_7 VPWR VGND sg13g2_decap_8
XFILLER_5_375 VPWR VGND sg13g2_decap_8
XFILLER_3_11 VPWR VGND sg13g2_decap_8
XFILLER_3_88 VPWR VGND sg13g2_decap_8
XFILLER_1_581 VPWR VGND sg13g2_decap_8
XFILLER_49_574 VPWR VGND sg13g2_decap_8
XFILLER_3_1028 VPWR VGND sg13g2_fill_1
XFILLER_36_268 VPWR VGND sg13g2_decap_8
XFILLER_37_769 VPWR VGND sg13g2_decap_8
XFILLER_33_964 VPWR VGND sg13g2_decap_8
XFILLER_20_614 VPWR VGND sg13g2_decap_8
XFILLER_32_474 VPWR VGND sg13g2_decap_8
XFILLER_47_28 VPWR VGND sg13g2_decap_8
XFILLER_27_224 VPWR VGND sg13g2_decap_8
XFILLER_28_736 VPWR VGND sg13g2_decap_8
XFILLER_16_909 VPWR VGND sg13g2_decap_8
XFILLER_24_942 VPWR VGND sg13g2_decap_8
XFILLER_23_452 VPWR VGND sg13g2_decap_8
XFILLER_10_102 VPWR VGND sg13g2_decap_8
XFILLER_11_669 VPWR VGND sg13g2_decap_8
X_080_ _034_ VPWR _047_ VGND _033_ mod1.i_out_8psk\[1\] sg13g2_o21ai_1
XFILLER_10_179 VPWR VGND sg13g2_decap_8
XFILLER_12_53 VPWR VGND sg13g2_decap_8
XFILLER_3_802 VPWR VGND sg13g2_decap_8
XFILLER_2_312 VPWR VGND sg13g2_decap_8
XFILLER_3_879 VPWR VGND sg13g2_decap_8
XFILLER_2_389 VPWR VGND sg13g2_decap_8
XFILLER_46_511 VPWR VGND sg13g2_decap_8
XFILLER_19_769 VPWR VGND sg13g2_decap_8
XFILLER_34_706 VPWR VGND sg13g2_decap_8
XFILLER_46_588 VPWR VGND sg13g2_decap_8
XFILLER_15_931 VPWR VGND sg13g2_decap_8
XFILLER_27_791 VPWR VGND sg13g2_decap_8
XFILLER_14_430 VPWR VGND sg13g2_decap_8
XFILLER_42_761 VPWR VGND sg13g2_decap_8
XFILLER_30_912 VPWR VGND sg13g2_decap_8
XFILLER_30_989 VPWR VGND sg13g2_decap_8
XFILLER_6_662 VPWR VGND sg13g2_decap_8
XFILLER_5_172 VPWR VGND sg13g2_decap_8
XFILLER_49_371 VPWR VGND sg13g2_decap_8
XFILLER_37_566 VPWR VGND sg13g2_decap_8
XFILLER_33_19 VPWR VGND sg13g2_decap_8
XFILLER_33_761 VPWR VGND sg13g2_decap_8
XFILLER_20_411 VPWR VGND sg13g2_decap_8
XFILLER_21_934 VPWR VGND sg13g2_decap_8
XFILLER_32_271 VPWR VGND sg13g2_decap_8
XFILLER_20_488 VPWR VGND sg13g2_decap_8
XFILLER_3_109 VPWR VGND sg13g2_decap_8
XFILLER_0_805 VPWR VGND sg13g2_decap_8
XFILLER_47_308 VPWR VGND sg13g2_decap_8
XFILLER_28_533 VPWR VGND sg13g2_decap_8
XFILLER_16_706 VPWR VGND sg13g2_decap_8
XFILLER_15_205 VPWR VGND sg13g2_decap_8
XFILLER_43_558 VPWR VGND sg13g2_decap_8
XFILLER_30_208 VPWR VGND sg13g2_decap_8
XFILLER_12_956 VPWR VGND sg13g2_decap_8
XFILLER_23_271 VPWR VGND sg13g2_decap_8
XFILLER_11_466 VPWR VGND sg13g2_decap_8
X_132_ net15 VGND VPWR mod1.qam16_mod.i_level\[3\] mod1.i_out_qam16\[3\] clknet_2_3__leaf_clk
+ sg13g2_dfrbpq_1
XFILLER_8_949 VPWR VGND sg13g2_decap_8
XFILLER_7_448 VPWR VGND sg13g2_decap_8
XFILLER_23_74 VPWR VGND sg13g2_decap_8
X_063_ net9 net8 _038_ VPWR VGND sg13g2_and2_1
XFILLER_3_676 VPWR VGND sg13g2_decap_8
XFILLER_2_186 VPWR VGND sg13g2_decap_8
XFILLER_39_809 VPWR VGND sg13g2_decap_8
XFILLER_38_319 VPWR VGND sg13g2_decap_8
XFILLER_47_875 VPWR VGND sg13g2_decap_8
XFILLER_19_566 VPWR VGND sg13g2_decap_8
XFILLER_46_385 VPWR VGND sg13g2_decap_8
XFILLER_0_56 VPWR VGND sg13g2_decap_8
XFILLER_34_503 VPWR VGND sg13g2_decap_8
XFILLER_22_709 VPWR VGND sg13g2_decap_8
XFILLER_9_32 VPWR VGND sg13g2_decap_8
XFILLER_30_786 VPWR VGND sg13g2_decap_8
XFILLER_9_1012 VPWR VGND sg13g2_decap_8
XFILLER_38_820 VPWR VGND sg13g2_decap_8
XFILLER_37_363 VPWR VGND sg13g2_fill_1
XFILLER_38_897 VPWR VGND sg13g2_decap_8
XFILLER_25_558 VPWR VGND sg13g2_decap_8
XFILLER_21_731 VPWR VGND sg13g2_decap_8
XFILLER_20_263 VPWR VGND sg13g2_decap_8
XFILLER_0_602 VPWR VGND sg13g2_decap_8
XFILLER_0_679 VPWR VGND sg13g2_decap_8
XFILLER_47_105 VPWR VGND sg13g2_decap_8
XFILLER_28_330 VPWR VGND sg13g2_fill_1
XFILLER_16_503 VPWR VGND sg13g2_decap_8
XFILLER_18_74 VPWR VGND sg13g2_decap_8
XFILLER_29_886 VPWR VGND sg13g2_decap_8
XFILLER_44_845 VPWR VGND sg13g2_decap_8
XFILLER_28_396 VPWR VGND sg13g2_decap_4
XFILLER_43_355 VPWR VGND sg13g2_decap_8
XFILLER_34_40 VPWR VGND sg13g2_decap_8
XFILLER_12_753 VPWR VGND sg13g2_decap_8
XFILLER_8_746 VPWR VGND sg13g2_decap_8
XFILLER_11_263 VPWR VGND sg13g2_decap_8
XFILLER_7_245 VPWR VGND sg13g2_decap_8
X_115_ net19 net18 net17 net1 _029_ VPWR VGND sg13g2_nor4_1
XFILLER_4_963 VPWR VGND sg13g2_decap_8
XFILLER_3_473 VPWR VGND sg13g2_decap_8
XFILLER_39_606 VPWR VGND sg13g2_decap_8
XFILLER_38_116 VPWR VGND sg13g2_decap_8
XFILLER_47_672 VPWR VGND sg13g2_decap_8
XFILLER_19_374 VPWR VGND sg13g2_decap_8
XFILLER_35_801 VPWR VGND sg13g2_decap_8
XFILLER_46_182 VPWR VGND sg13g2_decap_8
XFILLER_22_506 VPWR VGND sg13g2_decap_8
XFILLER_35_878 VPWR VGND sg13g2_decap_8
XFILLER_30_583 VPWR VGND sg13g2_decap_8
XFILLER_39_18 VPWR VGND sg13g2_decap_8
XFILLER_29_105 VPWR VGND sg13g2_decap_8
XFILLER_26_812 VPWR VGND sg13g2_decap_8
XFILLER_25_311 VPWR VGND sg13g2_decap_8
XFILLER_38_694 VPWR VGND sg13g2_decap_8
XFILLER_25_355 VPWR VGND sg13g2_fill_1
XFILLER_26_889 VPWR VGND sg13g2_decap_8
XFILLER_41_859 VPWR VGND sg13g2_decap_8
XFILLER_25_388 VPWR VGND sg13g2_decap_8
XFILLER_40_369 VPWR VGND sg13g2_decap_8
XFILLER_20_53 VPWR VGND sg13g2_decap_8
XFILLER_1_966 VPWR VGND sg13g2_decap_8
XFILLER_49_959 VPWR VGND sg13g2_decap_8
XFILLER_0_476 VPWR VGND sg13g2_decap_8
XFILLER_48_469 VPWR VGND sg13g2_decap_8
XFILLER_29_84 VPWR VGND sg13g2_decap_8
XFILLER_17_812 VPWR VGND sg13g2_decap_8
XFILLER_29_683 VPWR VGND sg13g2_decap_8
XFILLER_44_642 VPWR VGND sg13g2_decap_8
XFILLER_16_333 VPWR VGND sg13g2_decap_4
XFILLER_45_61 VPWR VGND sg13g2_decap_8
XFILLER_43_152 VPWR VGND sg13g2_decap_8
XFILLER_17_889 VPWR VGND sg13g2_decap_8
XFILLER_16_377 VPWR VGND sg13g2_decap_8
XFILLER_32_859 VPWR VGND sg13g2_decap_8
XFILLER_31_358 VPWR VGND sg13g2_decap_8
XFILLER_12_550 VPWR VGND sg13g2_decap_8
XFILLER_8_543 VPWR VGND sg13g2_decap_8
XFILLER_6_11 VPWR VGND sg13g2_decap_8
XFILLER_6_88 VPWR VGND sg13g2_decap_8
XFILLER_4_760 VPWR VGND sg13g2_decap_8
XFILLER_3_270 VPWR VGND sg13g2_decap_8
XFILLER_6_1026 VPWR VGND sg13g2_fill_2
XFILLER_39_403 VPWR VGND sg13g2_decap_8
XFILLER_27_609 VPWR VGND sg13g2_decap_8
XFILLER_34_152 VPWR VGND sg13g2_decap_8
XFILLER_35_675 VPWR VGND sg13g2_decap_8
XFILLER_23_837 VPWR VGND sg13g2_decap_8
XFILLER_22_369 VPWR VGND sg13g2_decap_8
XFILLER_30_380 VPWR VGND sg13g2_decap_8
Xheichips25_template_31 VPWR VGND uio_out[7] sg13g2_tielo
XFILLER_39_970 VPWR VGND sg13g2_decap_8
XFILLER_45_439 VPWR VGND sg13g2_decap_8
XFILLER_17_119 VPWR VGND sg13g2_decap_8
XFILLER_38_491 VPWR VGND sg13g2_decap_8
XFILLER_14_815 VPWR VGND sg13g2_decap_8
XFILLER_25_130 VPWR VGND sg13g2_decap_8
XFILLER_26_686 VPWR VGND sg13g2_decap_8
XFILLER_41_656 VPWR VGND sg13g2_decap_8
XFILLER_13_347 VPWR VGND sg13g2_decap_8
XFILLER_15_53 VPWR VGND sg13g2_decap_8
XFILLER_25_196 VPWR VGND sg13g2_decap_8
XFILLER_40_144 VPWR VGND sg13g2_decap_8
XFILLER_22_870 VPWR VGND sg13g2_decap_8
XFILLER_5_557 VPWR VGND sg13g2_decap_8
XFILLER_31_96 VPWR VGND sg13g2_decap_8
XFILLER_1_763 VPWR VGND sg13g2_decap_8
XFILLER_0_273 VPWR VGND sg13g2_decap_8
XFILLER_49_756 VPWR VGND sg13g2_decap_8
XFILLER_48_266 VPWR VGND sg13g2_decap_8
XFILLER_36_417 VPWR VGND sg13g2_decap_8
XFILLER_29_480 VPWR VGND sg13g2_decap_8
XFILLER_16_130 VPWR VGND sg13g2_decap_8
XFILLER_17_686 VPWR VGND sg13g2_decap_8
XFILLER_32_656 VPWR VGND sg13g2_decap_8
XFILLER_31_166 VPWR VGND sg13g2_decap_8
XFILLER_9_830 VPWR VGND sg13g2_decap_8
XFILLER_8_340 VPWR VGND sg13g2_decap_8
XFILLER_28_1016 VPWR VGND sg13g2_decap_8
XFILLER_28_1027 VPWR VGND sg13g2_fill_2
XFILLER_39_200 VPWR VGND sg13g2_decap_8
.ends

